
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_windowed_reg_M4_N4_F4_naddr4_nbit8 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_windowed_reg_M4_N4_F4_naddr4_nbit8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_reg_M4_N4_F4_naddr4_nbit8.all;

entity windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_add_0 is

   port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (4 downto 0);  CO : out std_logic);

end windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_add_0;

architecture SYN_rpl of windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1 : XOR2_X1 port map( A => A(4), B => carry_4_port, Z => SUM(4));
   U2 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);
   U3 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_reg_M4_N4_F4_naddr4_nbit8.all;

entity windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_2 is

   port( A, B : in std_logic_vector (5 downto 0);  CI, ADD_SUB : in std_logic; 
         SUM : out std_logic_vector (5 downto 0);  CO : out std_logic);

end windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_2;

architecture SYN_rpl of windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port,
      B_AS_3_port, B_AS_2_port, B_AS_1_port, B_AS_0_port, n_1007 : std_logic;

begin
   
   U1_5 : FA_X1 port map( A => A(5), B => ADD_SUB, CI => carry_5_port, CO => 
                           n_1007, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => ADD_SUB, CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U2 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U3 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U4 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_reg_M4_N4_F4_naddr4_nbit8.all;

entity windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in std_logic;
         SUM : out std_logic_vector (31 downto 0);  CO : out std_logic);

end windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_1;

architecture SYN_rpl of windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_0_port, 
      n_1042 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => ADD_SUB, CI => carry_31_port, CO =>
                           n_1042, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => ADD_SUB, CI => carry_30_port, CO =>
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => ADD_SUB, CI => carry_29_port, CO =>
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => ADD_SUB, CI => carry_28_port, CO =>
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => ADD_SUB, CI => carry_27_port, CO =>
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => ADD_SUB, CI => carry_26_port, CO =>
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => ADD_SUB, CI => carry_25_port, CO =>
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => ADD_SUB, CI => carry_24_port, CO =>
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => ADD_SUB, CI => carry_23_port, CO =>
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => ADD_SUB, CI => carry_22_port, CO =>
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => ADD_SUB, CI => carry_21_port, CO =>
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => ADD_SUB, CI => carry_20_port, CO =>
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => ADD_SUB, CI => carry_19_port, CO =>
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => ADD_SUB, CI => carry_18_port, CO =>
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => ADD_SUB, CI => carry_17_port, CO =>
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => ADD_SUB, CI => carry_16_port, CO =>
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => ADD_SUB, CI => carry_15_port, CO =>
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => ADD_SUB, CI => carry_14_port, CO =>
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => ADD_SUB, CI => carry_13_port, CO =>
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => ADD_SUB, CI => carry_12_port, CO =>
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => ADD_SUB, CI => carry_11_port, CO =>
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => ADD_SUB, CI => carry_10_port, CO =>
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => ADD_SUB, CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => ADD_SUB, CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => ADD_SUB, CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => ADD_SUB, CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => ADD_SUB, CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => ADD_SUB, CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => ADD_SUB, CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => ADD_SUB, CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => ADD_SUB, CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : INV_X1 port map( A => ADD_SUB, ZN => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_reg_M4_N4_F4_naddr4_nbit8.all;

entity windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_0 is

   port( A, B : in std_logic_vector (5 downto 0);  CI, ADD_SUB : in std_logic; 
         SUM : out std_logic_vector (5 downto 0);  CO : out std_logic);

end windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_0;

architecture SYN_rpl of windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_AS_4_port, 
      B_AS_3_port, B_AS_2_port, B_AS_1_port, B_AS_0_port : std_logic;

begin
   
   U1_3 : FA_X1 port map( A => A(3), B => B_AS_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B_AS_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B_AS_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B_AS_0_port, CI => ADD_SUB, CO => 
                           carry_1_port, S => SUM(0));
   U1 : XOR2_X1 port map( A => B_AS_4_port, B => carry_4_port, Z => SUM(4));
   U2 : XOR2_X1 port map( A => B(5), B => ADD_SUB, Z => B_AS_4_port);
   U3 : XOR2_X1 port map( A => B(3), B => ADD_SUB, Z => B_AS_3_port);
   U4 : XOR2_X1 port map( A => B(2), B => ADD_SUB, Z => B_AS_2_port);
   U5 : XOR2_X1 port map( A => B(1), B => ADD_SUB, Z => B_AS_1_port);
   U6 : XOR2_X1 port map( A => B(0), B => ADD_SUB, Z => B_AS_0_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_reg_M4_N4_F4_naddr4_nbit8.all;

entity windowed_reg_M4_N4_F4_naddr4_nbit8 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (3 downto 0);  DATAIN : in 
         std_logic_vector (7 downto 0);  OUT1, OUT2 : out std_logic_vector (7 
         downto 0);  CALL, RET : in std_logic;  FILL, SPILL : out std_logic;  
         DATA_FROM_MEM : in std_logic_vector (7 downto 0);  DATA_TO_MEM : out 
         std_logic_vector (7 downto 0));

end windowed_reg_M4_N4_F4_naddr4_nbit8;

architecture SYN_Behavioral of windowed_reg_M4_N4_F4_naddr4_nbit8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_add_0
      port( A, B : in std_logic_vector (4 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (4 downto 0);  CO : out std_logic);
   end component;
   
   component windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_2
      port( A, B : in std_logic_vector (5 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (5 downto 0);  CO : out 
            std_logic);
   end component;
   
   component windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_1
      port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (31 downto 0);  CO : out 
            std_logic);
   end component;
   
   component windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_0
      port( A, B : in std_logic_vector (5 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (5 downto 0);  CO : out 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, CWP_4_port, CWP_3_port, CWP_2_port, 
      CWP_1_port, CWP_0_port, counter_31_port, counter_30_port, counter_29_port
      , counter_28_port, counter_27_port, counter_26_port, counter_25_port, 
      counter_24_port, counter_23_port, counter_22_port, counter_21_port, 
      counter_20_port, counter_19_port, counter_18_port, counter_17_port, 
      counter_16_port, counter_15_port, counter_14_port, counter_13_port, 
      counter_12_port, counter_11_port, counter_10_port, counter_9_port, 
      counter_8_port, counter_7_port, counter_6_port, counter_5_port, 
      counter_4_port, counter_3_port, counter_2_port, counter_1_port, 
      counter_0_port, N107, N108, N109, N110, N111, N302, N303, N310, N311, 
      N312, N1191, N1193, N1195, N1197, N1199, N1201, N1203, N1205, N1207, 
      N1209, N1211, N1213, N1215, N1217, N1219, N1221, N1223, N1225, N1227, 
      N1229, N1231, N1233, N1235, N1237, N1239, N1241, N1243, N1245, N1247, 
      N1249, N1251, N1253, N1725, N1726, N1727, N1728, N1729, N1730, n8, n11, 
      n24, n28, U3_U3_Z_0, U3_U3_Z_1, U3_U3_Z_2, U3_U3_Z_3, U3_U3_Z_5, 
      U3_U4_Z_0, U3_U20_Z_0, U3_U21_Z_0, U3_U21_Z_1, U3_U21_Z_2, U3_U21_Z_3, 
      U3_U21_Z_4, U3_U21_Z_5, U3_U22_Z_0, U3_U22_Z_1, U3_U22_Z_2, U3_U22_Z_3, 
      U3_U23_Z_0, n1258, n1259, n1329, n1330, n1331, n1332, n1333, n1334, n1335
      , n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, 
      n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
      n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, 
      n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, 
      n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, 
      n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, 
      n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
      n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, 
      n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, 
      n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, 
      n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
      n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, 
      n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, 
      n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, 
      n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, 
      n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, 
      n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
      n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
      n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
      n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, 
      n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, 
      n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, 
      n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, 
      n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
      n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, 
      n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, 
      n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, 
      n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
      n1724, n1725_port, n1726_port, n1727_port, n1728_port, n1729_port, 
      n1730_port, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739
      , n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
      n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
      n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
      n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
      n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
      n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
      n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
      n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
      n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
      n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, 
      n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
      n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, 
      n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, 
      n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
      n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
      n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
      n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
      n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
      n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
      n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, 
      n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, 
      n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, 
      n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, 
      n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
      n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, 
      n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, 
      n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, 
      n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
      n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, 
      n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, 
      n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, 
      n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, 
      n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, 
      n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
      n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, 
      n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
      n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, 
      n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, 
      n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, 
      n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, 
      n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, 
      n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, 
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n8 <= '0';
   n11 <= '0';
   n24 <= '0';
   n28 <= '0';
   counter_reg_0_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           counter_0_port, QN => n3568);
   CANSAVE_reg : DFF_X1 port map( D => n1810, CK => CLK, Q => n_1049, QN => 
                           n2222);
   Storing_reg : DFF_X1 port map( D => n1809, CK => CLK, Q => n2189, QN => 
                           n3583);
   SWP_reg_4_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => n3585, QN => 
                           n2080);
   SWP_reg_0_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => n3589, QN => 
                           n2188);
   SWP_reg_1_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => n3588, QN => 
                           n2082);
   SWP_reg_2_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => n3587, QN => 
                           n2187);
   firstStoring_reg : DFF_X1 port map( D => n1804, CK => CLK, Q => n_1050, QN 
                           => n3581);
   SWP_reg_3_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => n3586, QN => 
                           n2081);
   CWP_reg_5_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => n2239, QN => 
                           n3590);
   CANRESTORE_reg : DFF_X1 port map( D => n1801, CK => CLK, Q => n_1051, QN => 
                           n3548);
   CWP_reg_3_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => CWP_3_port, QN
                           => n1813);
   CWP_reg_1_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => CWP_1_port, QN
                           => n1815);
   CWP_reg_0_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => CWP_0_port, QN
                           => n1816);
   CWP_reg_2_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => CWP_2_port, QN
                           => n1814);
   CWP_reg_4_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => CWP_4_port, QN
                           => n1812);
   GLOBAL_REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1795, CK => CLK, Q =>
                           n2231, QN => n3547);
   GLOBAL_REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1794, CK => CLK, Q =>
                           n2233, QN => n3546);
   GLOBAL_REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1793, CK => CLK, Q =>
                           n2235, QN => n3545);
   GLOBAL_REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1792, CK => CLK, Q =>
                           n2237, QN => n3544);
   GLOBAL_REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1791, CK => CLK, Q =>
                           n2238, QN => n3543);
   GLOBAL_REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1790, CK => CLK, Q =>
                           n2236, QN => n3542);
   GLOBAL_REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1789, CK => CLK, Q =>
                           n2234, QN => n3541);
   GLOBAL_REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1788, CK => CLK, Q =>
                           n2232, QN => n3540);
   GLOBAL_REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1787, CK => CLK, Q =>
                           n2240, QN => n3539);
   GLOBAL_REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1786, CK => CLK, Q =>
                           n2242, QN => n3538);
   GLOBAL_REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1785, CK => CLK, Q =>
                           n2244, QN => n3537);
   GLOBAL_REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q =>
                           n2246, QN => n3536);
   GLOBAL_REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q =>
                           n2247, QN => n3535);
   GLOBAL_REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1782, CK => CLK, Q =>
                           n2245, QN => n3534);
   GLOBAL_REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1781, CK => CLK, Q =>
                           n2243, QN => n3533);
   GLOBAL_REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1780, CK => CLK, Q =>
                           n2241, QN => n3532);
   GLOBAL_REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1779, CK => CLK, Q =>
                           n3531, QN => n2320);
   GLOBAL_REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1778, CK => CLK, Q =>
                           n3530, QN => n2321);
   GLOBAL_REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1777, CK => CLK, Q =>
                           n3529, QN => n2322);
   GLOBAL_REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1776, CK => CLK, Q =>
                           n3528, QN => n2323);
   GLOBAL_REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1775, CK => CLK, Q =>
                           n3527, QN => n2324);
   GLOBAL_REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1774, CK => CLK, Q =>
                           n3526, QN => n2325);
   GLOBAL_REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1773, CK => CLK, Q =>
                           n3525, QN => n2326);
   GLOBAL_REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1772, CK => CLK, Q =>
                           n3524, QN => n2327);
   GLOBAL_REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1771, CK => CLK, Q =>
                           n3523, QN => n2312);
   GLOBAL_REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1770, CK => CLK, Q =>
                           n3522, QN => n2313);
   GLOBAL_REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1769, CK => CLK, Q =>
                           n3521, QN => n2314);
   GLOBAL_REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1768, CK => CLK, Q =>
                           n3520, QN => n2315);
   GLOBAL_REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1767, CK => CLK, Q =>
                           n3519, QN => n2316);
   GLOBAL_REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1766, CK => CLK, Q =>
                           n3518, QN => n2317);
   GLOBAL_REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1765, CK => CLK, Q =>
                           n3517, QN => n2318);
   GLOBAL_REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1764, CK => CLK, Q =>
                           n3516, QN => n2319);
   counter_reg_30_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           counter_30_port, QN => n3553);
   counter_reg_1_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           counter_1_port, QN => n3573);
   counter_reg_2_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           counter_2_port, QN => n3554);
   counter_reg_3_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           counter_3_port, QN => n3559);
   counter_reg_4_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           counter_4_port, QN => n3558);
   counter_reg_5_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           counter_5_port, QN => n3557);
   counter_reg_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           counter_6_port, QN => n3564);
   counter_reg_7_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           counter_7_port, QN => n3563);
   counter_reg_8_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           counter_8_port, QN => n3562);
   counter_reg_9_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           counter_9_port, QN => n3561);
   counter_reg_10_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           counter_10_port, QN => n3567);
   counter_reg_11_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           counter_11_port, QN => n3566);
   counter_reg_12_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           counter_12_port, QN => n3565);
   counter_reg_13_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           counter_13_port, QN => n3572);
   counter_reg_14_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           counter_14_port, QN => n3571);
   counter_reg_15_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           counter_15_port, QN => n3570);
   counter_reg_16_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           counter_16_port, QN => n3569);
   counter_reg_17_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           counter_17_port, QN => n3576);
   counter_reg_18_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           counter_18_port, QN => n3575);
   counter_reg_19_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           counter_19_port, QN => n3574);
   counter_reg_20_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           counter_20_port, QN => n3580);
   counter_reg_21_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           counter_21_port, QN => n3579);
   counter_reg_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           counter_22_port, QN => n3578);
   counter_reg_23_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           counter_23_port, QN => n3577);
   counter_reg_24_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           counter_24_port, QN => n3552);
   counter_reg_25_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           counter_25_port, QN => n3551);
   counter_reg_26_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           counter_26_port, QN => n3550);
   counter_reg_27_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           counter_27_port, QN => n3549);
   counter_reg_28_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           counter_28_port, QN => n3556);
   counter_reg_29_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           counter_29_port, QN => n3555);
   counter_reg_31_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           counter_31_port, QN => n3560);
   SWP_reg_5_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => n3584, QN => 
                           n_1052);
   Restoring_reg : DFF_X1 port map( D => n1731, CK => CLK, Q => n_1053, QN => 
                           n3582);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1730_port, CK => CLK, Q => 
                           n3515, QN => n2256);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1729_port, CK => CLK, Q => 
                           n3514, QN => n2258);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1728_port, CK => CLK, Q => 
                           n3513, QN => n2260);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1727_port, CK => CLK, Q => 
                           n3512, QN => n2262);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1726_port, CK => CLK, Q => 
                           n3511, QN => n2263);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1725_port, CK => CLK, Q => 
                           n3510, QN => n2261);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => n3509,
                           QN => n2259);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => n3508,
                           QN => n2257);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => n3507,
                           QN => n2132);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => n3506,
                           QN => n2136);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => n3505,
                           QN => n2140);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => n3504,
                           QN => n2144);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => n3503,
                           QN => n2146);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => n3502,
                           QN => n2142);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => n3501,
                           QN => n2138);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => n3500,
                           QN => n2134);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => n3499,
                           QN => n2288);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => n3498,
                           QN => n2290);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => n3497,
                           QN => n2292);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => n3496,
                           QN => n2294);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => n3495,
                           QN => n2295);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => n3494,
                           QN => n2293);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => n3493,
                           QN => n2291);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => n3492,
                           QN => n2289);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => n3491,
                           QN => n2179);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => n3490,
                           QN => n2181);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => n3489,
                           QN => n2183);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => n3488,
                           QN => n2185);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => n3487,
                           QN => n2186);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => n3486,
                           QN => n2184);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => n3485,
                           QN => n2182);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => n3484,
                           QN => n2180);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => n3483,
                           QN => n_1054);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => n3482,
                           QN => n_1055);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => n3481,
                           QN => n_1056);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => n3480,
                           QN => n_1057);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => n3479,
                           QN => n_1058);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => n3478,
                           QN => n_1059);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => n3477,
                           QN => n_1060);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => n3476,
                           QN => n_1061);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => n3475,
                           QN => n_1062);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => n3474,
                           QN => n_1063);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => n3473,
                           QN => n_1064);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => n3472,
                           QN => n_1065);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => n3471,
                           QN => n_1066);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => n3470,
                           QN => n_1067);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => n3469,
                           QN => n_1068);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => n3468,
                           QN => n_1069);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => n3467,
                           QN => n2147);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => n3466,
                           QN => n2149);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => n3465,
                           QN => n2151);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => n3464,
                           QN => n2153);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => n3463,
                           QN => n2154);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => n3462,
                           QN => n2152);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => n3461,
                           QN => n2150);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => n3460,
                           QN => n2148);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => n3459,
                           QN => n2264);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => n3458,
                           QN => n2266);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => n3457,
                           QN => n2268);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => n3456,
                           QN => n2270);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => n3455,
                           QN => n2271);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => n3454,
                           QN => n2269);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => n3453,
                           QN => n2267);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => n3452,
                           QN => n2265);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => n3451,
                           QN => n2248);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => n3450,
                           QN => n2250);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => n3449,
                           QN => n2252);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => n3448,
                           QN => n2254);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => n3447,
                           QN => n2255);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => n3446,
                           QN => n2253);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => n3445,
                           QN => n2251);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => n3444,
                           QN => n2249);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => n3443,
                           QN => n2131);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => n3442,
                           QN => n2135);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => n3441,
                           QN => n2139);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => n3440,
                           QN => n2143);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => n3439,
                           QN => n2145);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => n3438,
                           QN => n2141);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => n3437,
                           QN => n2137);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => n3436,
                           QN => n2133);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => n3435
                           , QN => n2171);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => n3434
                           , QN => n2173);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => n3433
                           , QN => n2175);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => n3432
                           , QN => n2177);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => n3431
                           , QN => n2178);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => n3430
                           , QN => n2176);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => n3429
                           , QN => n2174);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => n3428
                           , QN => n2172);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => n3427
                           , QN => n2296);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => n3426
                           , QN => n2298);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => n3425
                           , QN => n2300);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => n3424
                           , QN => n2302);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => n3423
                           , QN => n2303);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => n3422
                           , QN => n2301);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => n3421
                           , QN => n2299);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => n3420
                           , QN => n2297);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => n3419
                           , QN => n_1070);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => n3418
                           , QN => n_1071);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => n3417
                           , QN => n_1072);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => n3416
                           , QN => n_1073);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => n3415
                           , QN => n_1074);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => n3414
                           , QN => n_1075);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n3413
                           , QN => n_1076);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => n3412
                           , QN => n_1077);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n3411
                           , QN => n_1078);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => n3410
                           , QN => n_1079);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n3409
                           , QN => n_1080);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => n3408
                           , QN => n_1081);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n3407
                           , QN => n_1082);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => n3406
                           , QN => n_1083);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n3405
                           , QN => n_1084);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => n3404
                           , QN => n_1085);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n3403
                           , QN => n2123);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => n3402
                           , QN => n2125);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n3401
                           , QN => n2127);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => n3400
                           , QN => n2129);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n3399
                           , QN => n2130);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => n3398
                           , QN => n2128);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n3397
                           , QN => n2126);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => n3396
                           , QN => n2124);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n3395
                           , QN => n2272);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => n3394
                           , QN => n2274);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n3393
                           , QN => n2276);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => n3392
                           , QN => n2278);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n3391
                           , QN => n2279);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => n3390
                           , QN => n2277);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n3389
                           , QN => n2275);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => n3388
                           , QN => n2273);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n3387
                           , QN => n2280);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => n3386
                           , QN => n2282);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n3385
                           , QN => n2284);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => n3384
                           , QN => n2286);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n3383
                           , QN => n2287);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => n3382
                           , QN => n2285);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n3381
                           , QN => n2283);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => n3380
                           , QN => n2281);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n3379
                           , QN => n2155);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => n3378
                           , QN => n2157);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n3377
                           , QN => n2159);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => n3376
                           , QN => n2161);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n3375
                           , QN => n2162);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => n3374
                           , QN => n2160);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n3373
                           , QN => n2158);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => n3372
                           , QN => n2156);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n3371
                           , QN => n2099);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => n3370
                           , QN => n2101);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n3369
                           , QN => n2103);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => n3368
                           , QN => n2105);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n3367
                           , QN => n2106);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => n3366
                           , QN => n2104);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n3365
                           , QN => n2102);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => n3364
                           , QN => n2100);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n3363
                           , QN => n2214);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => n3362
                           , QN => n2216);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n3361
                           , QN => n2218);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => n3360
                           , QN => n2220);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n3359
                           , QN => n2221);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => n3358
                           , QN => n2219);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n3357
                           , QN => n2217);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => n3356
                           , QN => n2215);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n3355
                           , QN => n2199);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => n3354
                           , QN => n2203);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n3353
                           , QN => n2207);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => n3352
                           , QN => n2211);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n3351
                           , QN => n2213);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => n3350
                           , QN => n2209);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n3349
                           , QN => n2205);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => n3348
                           , QN => n2201);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n3347
                           , QN => n2108);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => n3346
                           , QN => n2112);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n3345
                           , QN => n2116);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => n3344
                           , QN => n2120);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n3343
                           , QN => n2122);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => n3342
                           , QN => n2118);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n3341
                           , QN => n2114);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => n3340
                           , QN => n2110);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n3339
                           , QN => n_1086);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => n3338
                           , QN => n_1087);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n3337
                           , QN => n_1088);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => n3336
                           , QN => n_1089);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n3335
                           , QN => n_1090);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => n3334
                           , QN => n_1091);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n3333
                           , QN => n_1092);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => n3332
                           , QN => n_1093);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n3331
                           , QN => n_1094);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => n3330
                           , QN => n_1095);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n3329
                           , QN => n_1096);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => n3328
                           , QN => n_1097);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n3327
                           , QN => n_1098);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => n3326
                           , QN => n_1099);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n3325
                           , QN => n_1100);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => n3324
                           , QN => n_1101);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n3323
                           , QN => n2198);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => n3322
                           , QN => n2202);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n3321
                           , QN => n2206);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => n3320
                           , QN => n2210);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n3319
                           , QN => n2212);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => n3318
                           , QN => n2208);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n3317
                           , QN => n2204);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => n3316
                           , QN => n2200);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n3315
                           , QN => n2107);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => n3314
                           , QN => n2111);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n3313
                           , QN => n2115);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => n3312
                           , QN => n2119);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n3311
                           , QN => n2121);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => n3310
                           , QN => n2117);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n3309
                           , QN => n2113);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => n3308
                           , QN => n2109);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n3307
                           , QN => n2091);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => n3306
                           , QN => n2093);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n3305
                           , QN => n2095);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => n3304
                           , QN => n2097);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n3303
                           , QN => n2098);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => n3302
                           , QN => n2096);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n3301
                           , QN => n2094);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => n3300
                           , QN => n2092);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n3299
                           , QN => n2223);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => n3298
                           , QN => n2225);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n3297
                           , QN => n2227);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => n3296
                           , QN => n2229);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n3295
                           , QN => n2230);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => n3294
                           , QN => n2228);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n3293
                           , QN => n2226);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => n3292
                           , QN => n2224);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n3291
                           , QN => n2163);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => n3290
                           , QN => n2165);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n3289
                           , QN => n2167);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => n3288
                           , QN => n2169);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n3287
                           , QN => n2170);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n3286
                           , QN => n2168);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n3285
                           , QN => n2166);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n3284
                           , QN => n2164);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n3283
                           , QN => n2304);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n3282
                           , QN => n2306);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n3281
                           , QN => n2308);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n3280
                           , QN => n2310);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n3279
                           , QN => n2311);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n3278
                           , QN => n2309);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n3277
                           , QN => n2307);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n3276
                           , QN => n2305);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n2190
                           , QN => n_1102);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n2192
                           , QN => n_1103);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n2194
                           , QN => n_1104);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n2196
                           , QN => n_1105);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n2197
                           , QN => n_1106);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n2195
                           , QN => n_1107);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n2193
                           , QN => n_1108);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n2191
                           , QN => n_1109);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n2083
                           , QN => n_1110);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n2085
                           , QN => n_1111);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n2087
                           , QN => n_1112);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n2089
                           , QN => n_1113);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n2090
                           , QN => n_1114);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n2088
                           , QN => n_1115);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n2086
                           , QN => n_1116);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n2084
                           , QN => n_1117);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n1329, QN => 
                           n2352);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           n1330, QN => n2328);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n1331, QN => 
                           n2353);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           n1332, QN => n2329);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n1333, QN => 
                           n2354);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           n1334, QN => n2330);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n1335, QN => 
                           n2355);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           n1336, QN => n2331);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n1337, QN => 
                           n2356);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           n1338, QN => n2332);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n1339, QN => 
                           n2357);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           n1340, QN => n2333);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n1341, QN => 
                           n2358);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           n1342, QN => n2334);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n1343, QN => 
                           n2359);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           n1344, QN => n2335);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n1345, QN => 
                           n2360);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           n1346, QN => n2336);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n1347, QN => 
                           n2361);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           n1348, QN => n2337);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n1349, QN => 
                           n2362);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           n1350, QN => n2338);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n1351, QN => 
                           n2363);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           n1352, QN => n2339);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n1353, QN => 
                           n2364);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           n1354, QN => n2340);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n1355, QN => 
                           n2365);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           n1356, QN => n2341);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n1357, QN => 
                           n2366);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           n1358, QN => n2342);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n1359, QN => 
                           n2367);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           n1360, QN => n2343);
   DATA_TO_MEM_reg_7_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n1361,
                           QN => n_1118);
   DATA_TO_MEM_tri_enable_reg_7_inst : DFF_X1 port map( D => n1441, CK => CLK, 
                           Q => n1362, QN => n2344);
   DATA_TO_MEM_reg_6_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n1363,
                           QN => n_1119);
   DATA_TO_MEM_tri_enable_reg_6_inst : DFF_X1 port map( D => n1439, CK => CLK, 
                           Q => n1364, QN => n2345);
   DATA_TO_MEM_reg_5_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n1365,
                           QN => n_1120);
   DATA_TO_MEM_tri_enable_reg_5_inst : DFF_X1 port map( D => n1437, CK => CLK, 
                           Q => n1366, QN => n2346);
   DATA_TO_MEM_reg_4_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n1367,
                           QN => n_1121);
   DATA_TO_MEM_tri_enable_reg_4_inst : DFF_X1 port map( D => n1435, CK => CLK, 
                           Q => n1368, QN => n2347);
   DATA_TO_MEM_reg_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n1369,
                           QN => n_1122);
   DATA_TO_MEM_tri_enable_reg_3_inst : DFF_X1 port map( D => n1433, CK => CLK, 
                           Q => n1370, QN => n2348);
   DATA_TO_MEM_reg_2_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n1371,
                           QN => n_1123);
   DATA_TO_MEM_tri_enable_reg_2_inst : DFF_X1 port map( D => n1431, CK => CLK, 
                           Q => n1372, QN => n2349);
   DATA_TO_MEM_reg_1_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n1373,
                           QN => n_1124);
   DATA_TO_MEM_tri_enable_reg_1_inst : DFF_X1 port map( D => n1429, CK => CLK, 
                           Q => n1374, QN => n2350);
   DATA_TO_MEM_reg_0_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n1375,
                           QN => n_1125);
   DATA_TO_MEM_tri_enable_reg_0_inst : DFF_X1 port map( D => n1427, CK => CLK, 
                           Q => n1376, QN => n2351);
   FILL_reg : DFF_X1 port map( D => n1426, CK => CLK, Q => FILL, QN => n1259);
   SPILL_reg : DFF_X1 port map( D => n1425, CK => CLK, Q => SPILL, QN => n1258)
                           ;
   r189 : windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_0 port map( A(5) => 
                           X_Logic0_port, A(4) => X_Logic0_port, A(3) => 
                           ADD_WR(3), A(2) => ADD_WR(2), A(1) => ADD_WR(1), 
                           A(0) => ADD_WR(0), B(5) => U3_U3_Z_5, B(4) => 
                           U3_U3_Z_5, B(3) => U3_U3_Z_3, B(2) => U3_U3_Z_2, 
                           B(1) => U3_U3_Z_1, B(0) => U3_U3_Z_0, CI => n8, 
                           ADD_SUB => U3_U4_Z_0, SUM(5) => n_1126, SUM(4) => 
                           N312, SUM(3) => N311, SUM(2) => N310, SUM(1) => N303
                           , SUM(0) => N302, CO => n_1127);
   r198 : windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_1 port map( A(31) => 
                           counter_31_port, A(30) => counter_30_port, A(29) => 
                           counter_29_port, A(28) => counter_28_port, A(27) => 
                           counter_27_port, A(26) => counter_26_port, A(25) => 
                           counter_25_port, A(24) => counter_24_port, A(23) => 
                           counter_23_port, A(22) => counter_22_port, A(21) => 
                           counter_21_port, A(20) => counter_20_port, A(19) => 
                           counter_19_port, A(18) => counter_18_port, A(17) => 
                           counter_17_port, A(16) => counter_16_port, A(15) => 
                           counter_15_port, A(14) => counter_14_port, A(13) => 
                           counter_13_port, A(12) => counter_12_port, A(11) => 
                           counter_11_port, A(10) => counter_10_port, A(9) => 
                           counter_9_port, A(8) => counter_8_port, A(7) => 
                           counter_7_port, A(6) => counter_6_port, A(5) => 
                           counter_5_port, A(4) => counter_4_port, A(3) => 
                           counter_3_port, A(2) => counter_2_port, A(1) => 
                           counter_1_port, A(0) => counter_0_port, B(31) => 
                           X_Logic0_port, B(30) => X_Logic0_port, B(29) => 
                           X_Logic0_port, B(28) => X_Logic0_port, B(27) => 
                           X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
                           X_Logic0_port, B(24) => X_Logic0_port, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic1_port, CI => n11, 
                           ADD_SUB => U3_U20_Z_0, SUM(31) => N1253, SUM(30) => 
                           N1251, SUM(29) => N1249, SUM(28) => N1247, SUM(27) 
                           => N1245, SUM(26) => N1243, SUM(25) => N1241, 
                           SUM(24) => N1239, SUM(23) => N1237, SUM(22) => N1235
                           , SUM(21) => N1233, SUM(20) => N1231, SUM(19) => 
                           N1229, SUM(18) => N1227, SUM(17) => N1225, SUM(16) 
                           => N1223, SUM(15) => N1221, SUM(14) => N1219, 
                           SUM(13) => N1217, SUM(12) => N1215, SUM(11) => N1213
                           , SUM(10) => N1211, SUM(9) => N1209, SUM(8) => N1207
                           , SUM(7) => N1205, SUM(6) => N1203, SUM(5) => N1201,
                           SUM(4) => N1199, SUM(3) => N1197, SUM(2) => N1195, 
                           SUM(1) => N1193, SUM(0) => N1191, CO => n_1128);
   r197 : windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_addsub_2 port map( A(5) => 
                           U3_U21_Z_5, A(4) => U3_U21_Z_4, A(3) => U3_U21_Z_3, 
                           A(2) => U3_U21_Z_2, A(1) => U3_U21_Z_1, A(0) => 
                           U3_U21_Z_0, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => U3_U22_Z_3, B(2) => 
                           U3_U22_Z_2, B(1) => U3_U22_Z_1, B(0) => U3_U22_Z_0, 
                           CI => n24, ADD_SUB => U3_U23_Z_0, SUM(5) => N1730, 
                           SUM(4) => N1729, SUM(3) => N1728, SUM(2) => N1727, 
                           SUM(1) => N1726, SUM(0) => N1725, CO => n_1129);
   add_168 : windowed_reg_M4_N4_F4_naddr4_nbit8_DW01_add_0 port map( A(4) => 
                           CWP_4_port, A(3) => CWP_3_port, A(2) => CWP_2_port, 
                           A(1) => CWP_1_port, A(0) => CWP_0_port, B(4) => 
                           X_Logic0_port, B(3) => ADD_RD1(3), B(2) => 
                           ADD_RD1(2), B(1) => ADD_RD1(1), B(0) => ADD_RD1(0), 
                           CI => n28, SUM(4) => N111, SUM(3) => N110, SUM(2) =>
                           N109, SUM(1) => N108, SUM(0) => N107, CO => n_1130);
   DATA_TO_MEM_tri_0_inst : TBUF_X1 port map( A => n1375, EN => n1376, Z => 
                           DATA_TO_MEM(0));
   DATA_TO_MEM_tri_1_inst : TBUF_X1 port map( A => n1373, EN => n1374, Z => 
                           DATA_TO_MEM(1));
   DATA_TO_MEM_tri_2_inst : TBUF_X1 port map( A => n1371, EN => n1372, Z => 
                           DATA_TO_MEM(2));
   DATA_TO_MEM_tri_3_inst : TBUF_X1 port map( A => n1369, EN => n1370, Z => 
                           DATA_TO_MEM(3));
   DATA_TO_MEM_tri_4_inst : TBUF_X1 port map( A => n1367, EN => n1368, Z => 
                           DATA_TO_MEM(4));
   DATA_TO_MEM_tri_5_inst : TBUF_X1 port map( A => n1365, EN => n1366, Z => 
                           DATA_TO_MEM(5));
   DATA_TO_MEM_tri_6_inst : TBUF_X1 port map( A => n1363, EN => n1364, Z => 
                           DATA_TO_MEM(6));
   DATA_TO_MEM_tri_7_inst : TBUF_X1 port map( A => n1361, EN => n1362, Z => 
                           DATA_TO_MEM(7));
   OUT2_tri_0_inst : TBUF_X1 port map( A => n1359, EN => n1360, Z => OUT2(0));
   OUT2_tri_1_inst : TBUF_X1 port map( A => n1357, EN => n1358, Z => OUT2(1));
   OUT2_tri_2_inst : TBUF_X1 port map( A => n1355, EN => n1356, Z => OUT2(2));
   OUT2_tri_3_inst : TBUF_X1 port map( A => n1353, EN => n1354, Z => OUT2(3));
   OUT2_tri_4_inst : TBUF_X1 port map( A => n1351, EN => n1352, Z => OUT2(4));
   OUT2_tri_5_inst : TBUF_X1 port map( A => n1349, EN => n1350, Z => OUT2(5));
   OUT2_tri_6_inst : TBUF_X1 port map( A => n1347, EN => n1348, Z => OUT2(6));
   OUT2_tri_7_inst : TBUF_X1 port map( A => n1345, EN => n1346, Z => OUT2(7));
   OUT1_tri_0_inst : TBUF_X1 port map( A => n1343, EN => n1344, Z => OUT1(0));
   OUT1_tri_1_inst : TBUF_X1 port map( A => n1341, EN => n1342, Z => OUT1(1));
   OUT1_tri_2_inst : TBUF_X1 port map( A => n1339, EN => n1340, Z => OUT1(2));
   OUT1_tri_3_inst : TBUF_X1 port map( A => n1337, EN => n1338, Z => OUT1(3));
   OUT1_tri_4_inst : TBUF_X1 port map( A => n1335, EN => n1336, Z => OUT1(4));
   OUT1_tri_5_inst : TBUF_X1 port map( A => n1333, EN => n1334, Z => OUT1(5));
   OUT1_tri_6_inst : TBUF_X1 port map( A => n1331, EN => n1332, Z => OUT1(6));
   OUT1_tri_7_inst : TBUF_X1 port map( A => n1329, EN => n1330, Z => OUT1(7));
   U1676 : NAND2_X2 port map( A1 => n2374, A2 => n2368, ZN => n2369);
   U1677 : NAND3_X2 port map( A1 => n2464, A2 => n2374, A3 => n2465, ZN => 
                           n2368);
   U1678 : NAND2_X4 port map( A1 => CALL, A2 => n3275, ZN => U3_U20_Z_0);
   U1679 : INV_X4 port map( A => RESET, ZN => n2374);
   U1680 : OAI22_X1 port map( A1 => n3568, A2 => n2368, B1 => n2369, B2 => 
                           n2370, ZN => n1811);
   U1681 : INV_X1 port map( A => N1191, ZN => n2370);
   U1682 : OAI221_X1 port map( B1 => n2371, B2 => n2372, C1 => n2373, C2 => 
                           n2222, A => n2374, ZN => n1810);
   U1683 : NOR4_X1 port map( A1 => n1812, A2 => n2375, A3 => n2376, A4 => 
                           CWP_3_port, ZN => n2373);
   U1684 : OAI21_X1 port map( B1 => n3583, B2 => n2377, A => n2378, ZN => n1809
                           );
   U1685 : OAI221_X1 port map( B1 => n2379, B2 => n2380, C1 => n2381, C2 => 
                           n2080, A => n2382, ZN => n1808);
   U1686 : OAI221_X1 port map( B1 => n2379, B2 => n2383, C1 => n2381, C2 => 
                           n2188, A => n2382, ZN => n1807);
   U1687 : OAI221_X1 port map( B1 => n2379, B2 => n2384, C1 => n2381, C2 => 
                           n2082, A => n2382, ZN => n1806);
   U1688 : OAI221_X1 port map( B1 => n2379, B2 => n2385, C1 => n2381, C2 => 
                           n2187, A => n2382, ZN => n1805);
   U1689 : NAND2_X1 port map( A1 => n2386, A2 => n2374, ZN => n1804);
   U1690 : MUX2_X1 port map( A => n3581, B => n2387, S => n2388, Z => n2386);
   U1691 : NOR2_X1 port map( A1 => n2389, A2 => n2390, ZN => n2388);
   U1692 : OAI221_X1 port map( B1 => n2379, B2 => n2391, C1 => n2381, C2 => 
                           n2081, A => n2382, ZN => n1803);
   U1693 : NAND3_X1 port map( A1 => n2392, A2 => n3583, A3 => n2393, ZN => 
                           n2382);
   U1694 : INV_X1 port map( A => n2393, ZN => n2379);
   U1695 : OAI21_X1 port map( B1 => n3590, B2 => n2394, A => n2395, ZN => n1802
                           );
   U1696 : NAND4_X1 port map( A1 => N1730, A2 => n2396, A3 => U3_U20_Z_0, A4 =>
                           n2397, ZN => n2395);
   U1697 : AOI211_X1 port map( C1 => n3548, C2 => n2376, A => RESET, B => n2398
                           , ZN => n1801);
   U1698 : NOR3_X1 port map( A1 => n2399, A2 => CALL, A3 => n2400, ZN => n2398)
                           ;
   U1699 : OAI21_X1 port map( B1 => n1813, B2 => n2394, A => n2401, ZN => n1800
                           );
   U1700 : OAI21_X1 port map( B1 => n2402, B2 => N1728, A => n2396, ZN => n2401
                           );
   U1701 : OAI22_X1 port map( A1 => n1815, A2 => n2394, B1 => n2384, B2 => 
                           n2403, ZN => n1799);
   U1702 : OAI22_X1 port map( A1 => n1816, A2 => n2394, B1 => n2383, B2 => 
                           n2403, ZN => n1798);
   U1703 : OAI22_X1 port map( A1 => n1814, A2 => n2394, B1 => n2385, B2 => 
                           n2403, ZN => n1797);
   U1704 : NAND2_X1 port map( A1 => n2396, A2 => n2404, ZN => n2403);
   U1705 : OAI21_X1 port map( B1 => n1812, B2 => n2394, A => n2405, ZN => n1796
                           );
   U1706 : OAI21_X1 port map( B1 => n2402, B2 => N1729, A => n2396, ZN => n2405
                           );
   U1707 : AND2_X1 port map( A1 => n2374, A2 => n2394, ZN => n2396);
   U1708 : INV_X1 port map( A => n2404, ZN => n2402);
   U1709 : NAND2_X1 port map( A1 => n2406, A2 => U3_U20_Z_0, ZN => n2404);
   U1710 : OAI211_X1 port map( C1 => n2407, C2 => n2371, A => n2376, B => n2374
                           , ZN => n2394);
   U1711 : INV_X1 port map( A => n2408, ZN => n2371);
   U1712 : OAI22_X1 port map( A1 => n3547, A2 => n2409, B1 => n2410, B2 => 
                           n2411, ZN => n1795);
   U1713 : OAI22_X1 port map( A1 => n3546, A2 => n2409, B1 => n2410, B2 => 
                           n2412, ZN => n1794);
   U1714 : OAI22_X1 port map( A1 => n3545, A2 => n2409, B1 => n2410, B2 => 
                           n2413, ZN => n1793);
   U1715 : OAI22_X1 port map( A1 => n3544, A2 => n2409, B1 => n2410, B2 => 
                           n2414, ZN => n1792);
   U1716 : OAI22_X1 port map( A1 => n3543, A2 => n2409, B1 => n2410, B2 => 
                           n2415, ZN => n1791);
   U1717 : OAI22_X1 port map( A1 => n3542, A2 => n2409, B1 => n2410, B2 => 
                           n2416, ZN => n1790);
   U1718 : OAI22_X1 port map( A1 => n3541, A2 => n2409, B1 => n2410, B2 => 
                           n2417, ZN => n1789);
   U1719 : OAI22_X1 port map( A1 => n3540, A2 => n2409, B1 => n2410, B2 => 
                           n2418, ZN => n1788);
   U1720 : NAND2_X1 port map( A1 => n2374, A2 => n2409, ZN => n2410);
   U1721 : NAND2_X1 port map( A1 => n2374, A2 => n2419, ZN => n2409);
   U1722 : NAND3_X1 port map( A1 => n2420, A2 => n2421, A3 => n2422, ZN => 
                           n2419);
   U1723 : OAI22_X1 port map( A1 => n3539, A2 => n2423, B1 => n2411, B2 => 
                           n2424, ZN => n1787);
   U1724 : OAI22_X1 port map( A1 => n3538, A2 => n2423, B1 => n2412, B2 => 
                           n2424, ZN => n1786);
   U1725 : OAI22_X1 port map( A1 => n3537, A2 => n2423, B1 => n2413, B2 => 
                           n2424, ZN => n1785);
   U1726 : OAI22_X1 port map( A1 => n3536, A2 => n2423, B1 => n2414, B2 => 
                           n2424, ZN => n1784);
   U1727 : OAI22_X1 port map( A1 => n3535, A2 => n2423, B1 => n2415, B2 => 
                           n2424, ZN => n1783);
   U1728 : OAI22_X1 port map( A1 => n3534, A2 => n2423, B1 => n2416, B2 => 
                           n2424, ZN => n1782);
   U1729 : OAI22_X1 port map( A1 => n3533, A2 => n2423, B1 => n2417, B2 => 
                           n2424, ZN => n1781);
   U1730 : OAI22_X1 port map( A1 => n3532, A2 => n2423, B1 => n2418, B2 => 
                           n2424, ZN => n1780);
   U1731 : NAND2_X1 port map( A1 => n2374, A2 => n2423, ZN => n2424);
   U1732 : NAND2_X1 port map( A1 => n2374, A2 => n2425, ZN => n2423);
   U1733 : NAND3_X1 port map( A1 => n2422, A2 => n2421, A3 => N302, ZN => n2425
                           );
   U1734 : OAI22_X1 port map( A1 => n2426, A2 => n2320, B1 => n2411, B2 => 
                           n2427, ZN => n1779);
   U1735 : OAI22_X1 port map( A1 => n2426, A2 => n2321, B1 => n2412, B2 => 
                           n2427, ZN => n1778);
   U1736 : OAI22_X1 port map( A1 => n2426, A2 => n2322, B1 => n2413, B2 => 
                           n2427, ZN => n1777);
   U1737 : OAI22_X1 port map( A1 => n2426, A2 => n2323, B1 => n2414, B2 => 
                           n2427, ZN => n1776);
   U1738 : OAI22_X1 port map( A1 => n2426, A2 => n2324, B1 => n2415, B2 => 
                           n2427, ZN => n1775);
   U1739 : OAI22_X1 port map( A1 => n2426, A2 => n2325, B1 => n2416, B2 => 
                           n2427, ZN => n1774);
   U1740 : OAI22_X1 port map( A1 => n2426, A2 => n2326, B1 => n2417, B2 => 
                           n2427, ZN => n1773);
   U1741 : OAI22_X1 port map( A1 => n2426, A2 => n2327, B1 => n2418, B2 => 
                           n2427, ZN => n1772);
   U1742 : NAND2_X1 port map( A1 => n2374, A2 => n2426, ZN => n2427);
   U1743 : NAND2_X1 port map( A1 => n2374, A2 => n2428, ZN => n2426);
   U1744 : NAND3_X1 port map( A1 => n2422, A2 => n2420, A3 => N303, ZN => n2428
                           );
   U1745 : OAI22_X1 port map( A1 => n2429, A2 => n2312, B1 => n2411, B2 => 
                           n2430, ZN => n1771);
   U1746 : INV_X1 port map( A => DATAIN(7), ZN => n2411);
   U1747 : OAI22_X1 port map( A1 => n2429, A2 => n2313, B1 => n2412, B2 => 
                           n2430, ZN => n1770);
   U1748 : INV_X1 port map( A => DATAIN(5), ZN => n2412);
   U1749 : OAI22_X1 port map( A1 => n2429, A2 => n2314, B1 => n2413, B2 => 
                           n2430, ZN => n1769);
   U1750 : INV_X1 port map( A => DATAIN(3), ZN => n2413);
   U1751 : OAI22_X1 port map( A1 => n2429, A2 => n2315, B1 => n2414, B2 => 
                           n2430, ZN => n1768);
   U1752 : INV_X1 port map( A => DATAIN(1), ZN => n2414);
   U1753 : OAI22_X1 port map( A1 => n2429, A2 => n2316, B1 => n2415, B2 => 
                           n2430, ZN => n1767);
   U1754 : INV_X1 port map( A => DATAIN(0), ZN => n2415);
   U1755 : OAI22_X1 port map( A1 => n2429, A2 => n2317, B1 => n2416, B2 => 
                           n2430, ZN => n1766);
   U1756 : INV_X1 port map( A => DATAIN(2), ZN => n2416);
   U1757 : OAI22_X1 port map( A1 => n2429, A2 => n2318, B1 => n2417, B2 => 
                           n2430, ZN => n1765);
   U1758 : INV_X1 port map( A => DATAIN(4), ZN => n2417);
   U1759 : OAI22_X1 port map( A1 => n2429, A2 => n2319, B1 => n2418, B2 => 
                           n2430, ZN => n1764);
   U1760 : NAND2_X1 port map( A1 => n2374, A2 => n2429, ZN => n2430);
   U1761 : INV_X1 port map( A => DATAIN(6), ZN => n2418);
   U1762 : NAND2_X1 port map( A1 => n2374, A2 => n2431, ZN => n2429);
   U1763 : NAND3_X1 port map( A1 => N302, A2 => n2422, A3 => N303, ZN => n2431)
                           ;
   U1764 : AND3_X1 port map( A1 => U3_U4_Z_0, A2 => n2432, A3 => WR, ZN => 
                           n2422);
   U1765 : OAI22_X1 port map( A1 => n3553, A2 => n2368, B1 => n2369, B2 => 
                           n2433, ZN => n1763);
   U1766 : INV_X1 port map( A => N1251, ZN => n2433);
   U1767 : OAI22_X1 port map( A1 => n3573, A2 => n2368, B1 => n2369, B2 => 
                           n2434, ZN => n1762);
   U1768 : INV_X1 port map( A => N1193, ZN => n2434);
   U1769 : OAI22_X1 port map( A1 => n3554, A2 => n2368, B1 => n2369, B2 => 
                           n2435, ZN => n1761);
   U1770 : INV_X1 port map( A => N1195, ZN => n2435);
   U1771 : OAI22_X1 port map( A1 => n3559, A2 => n2368, B1 => n2369, B2 => 
                           n2436, ZN => n1760);
   U1772 : INV_X1 port map( A => N1197, ZN => n2436);
   U1773 : OAI22_X1 port map( A1 => n3558, A2 => n2368, B1 => n2369, B2 => 
                           n2437, ZN => n1759);
   U1774 : INV_X1 port map( A => N1199, ZN => n2437);
   U1775 : OAI22_X1 port map( A1 => n3557, A2 => n2368, B1 => n2369, B2 => 
                           n2438, ZN => n1758);
   U1776 : INV_X1 port map( A => N1201, ZN => n2438);
   U1777 : OAI22_X1 port map( A1 => n3564, A2 => n2368, B1 => n2369, B2 => 
                           n2439, ZN => n1757);
   U1778 : INV_X1 port map( A => N1203, ZN => n2439);
   U1779 : OAI22_X1 port map( A1 => n3563, A2 => n2368, B1 => n2369, B2 => 
                           n2440, ZN => n1756);
   U1780 : INV_X1 port map( A => N1205, ZN => n2440);
   U1781 : OAI22_X1 port map( A1 => n3562, A2 => n2368, B1 => n2369, B2 => 
                           n2441, ZN => n1755);
   U1782 : INV_X1 port map( A => N1207, ZN => n2441);
   U1783 : OAI22_X1 port map( A1 => n3561, A2 => n2368, B1 => n2369, B2 => 
                           n2442, ZN => n1754);
   U1784 : INV_X1 port map( A => N1209, ZN => n2442);
   U1785 : OAI22_X1 port map( A1 => n3567, A2 => n2368, B1 => n2369, B2 => 
                           n2443, ZN => n1753);
   U1786 : INV_X1 port map( A => N1211, ZN => n2443);
   U1787 : OAI22_X1 port map( A1 => n3566, A2 => n2368, B1 => n2369, B2 => 
                           n2444, ZN => n1752);
   U1788 : INV_X1 port map( A => N1213, ZN => n2444);
   U1789 : OAI22_X1 port map( A1 => n3565, A2 => n2368, B1 => n2369, B2 => 
                           n2445, ZN => n1751);
   U1790 : INV_X1 port map( A => N1215, ZN => n2445);
   U1791 : OAI22_X1 port map( A1 => n3572, A2 => n2368, B1 => n2369, B2 => 
                           n2446, ZN => n1750);
   U1792 : INV_X1 port map( A => N1217, ZN => n2446);
   U1793 : OAI22_X1 port map( A1 => n3571, A2 => n2368, B1 => n2369, B2 => 
                           n2447, ZN => n1749);
   U1794 : INV_X1 port map( A => N1219, ZN => n2447);
   U1795 : OAI22_X1 port map( A1 => n3570, A2 => n2368, B1 => n2369, B2 => 
                           n2448, ZN => n1748);
   U1796 : INV_X1 port map( A => N1221, ZN => n2448);
   U1797 : OAI22_X1 port map( A1 => n3569, A2 => n2368, B1 => n2369, B2 => 
                           n2449, ZN => n1747);
   U1798 : INV_X1 port map( A => N1223, ZN => n2449);
   U1799 : OAI22_X1 port map( A1 => n3576, A2 => n2368, B1 => n2369, B2 => 
                           n2450, ZN => n1746);
   U1800 : INV_X1 port map( A => N1225, ZN => n2450);
   U1801 : OAI22_X1 port map( A1 => n3575, A2 => n2368, B1 => n2369, B2 => 
                           n2451, ZN => n1745);
   U1802 : INV_X1 port map( A => N1227, ZN => n2451);
   U1803 : OAI22_X1 port map( A1 => n3574, A2 => n2368, B1 => n2369, B2 => 
                           n2452, ZN => n1744);
   U1804 : INV_X1 port map( A => N1229, ZN => n2452);
   U1805 : OAI22_X1 port map( A1 => n3580, A2 => n2368, B1 => n2369, B2 => 
                           n2453, ZN => n1743);
   U1806 : INV_X1 port map( A => N1231, ZN => n2453);
   U1807 : OAI22_X1 port map( A1 => n3579, A2 => n2368, B1 => n2369, B2 => 
                           n2454, ZN => n1742);
   U1808 : INV_X1 port map( A => N1233, ZN => n2454);
   U1809 : OAI22_X1 port map( A1 => n3578, A2 => n2368, B1 => n2369, B2 => 
                           n2455, ZN => n1741);
   U1810 : INV_X1 port map( A => N1235, ZN => n2455);
   U1811 : OAI22_X1 port map( A1 => n3577, A2 => n2368, B1 => n2369, B2 => 
                           n2456, ZN => n1740);
   U1812 : INV_X1 port map( A => N1237, ZN => n2456);
   U1813 : OAI22_X1 port map( A1 => n3552, A2 => n2368, B1 => n2369, B2 => 
                           n2457, ZN => n1739);
   U1814 : INV_X1 port map( A => N1239, ZN => n2457);
   U1815 : OAI22_X1 port map( A1 => n3551, A2 => n2368, B1 => n2369, B2 => 
                           n2458, ZN => n1738);
   U1816 : INV_X1 port map( A => N1241, ZN => n2458);
   U1817 : OAI22_X1 port map( A1 => n3550, A2 => n2368, B1 => n2369, B2 => 
                           n2459, ZN => n1737);
   U1818 : INV_X1 port map( A => N1243, ZN => n2459);
   U1819 : OAI22_X1 port map( A1 => n3549, A2 => n2368, B1 => n2369, B2 => 
                           n2460, ZN => n1736);
   U1820 : INV_X1 port map( A => N1245, ZN => n2460);
   U1821 : OAI22_X1 port map( A1 => n3556, A2 => n2368, B1 => n2369, B2 => 
                           n2461, ZN => n1735);
   U1822 : INV_X1 port map( A => N1247, ZN => n2461);
   U1823 : OAI22_X1 port map( A1 => n3555, A2 => n2368, B1 => n2369, B2 => 
                           n2462, ZN => n1734);
   U1824 : INV_X1 port map( A => N1249, ZN => n2462);
   U1825 : OAI22_X1 port map( A1 => n3560, A2 => n2368, B1 => n2369, B2 => 
                           n2463, ZN => n1733);
   U1826 : INV_X1 port map( A => N1253, ZN => n2463);
   U1827 : NAND3_X1 port map( A1 => n2406, A2 => n2372, A3 => n2408, ZN => 
                           n2465);
   U1828 : OR4_X1 port map( A1 => n2376, A2 => n2375, A3 => n1812, A4 => n1813,
                           ZN => n2464);
   U1829 : INV_X1 port map( A => n2466, ZN => n2376);
   U1830 : AOI21_X1 port map( B1 => n2467, B2 => n2468, A => n2392, ZN => n1732
                           );
   U1831 : NAND3_X1 port map( A1 => n2393, A2 => n3583, A3 => N1730, ZN => 
                           n2468);
   U1832 : NOR2_X1 port map( A1 => RESET, A2 => n2469, ZN => n2393);
   U1833 : NAND2_X1 port map( A1 => n3584, A2 => n2469, ZN => n2467);
   U1834 : INV_X1 port map( A => n2381, ZN => n2469);
   U1835 : OAI21_X1 port map( B1 => n2470, B2 => n2471, A => n2472, ZN => n2381
                           );
   U1836 : NOR2_X1 port map( A1 => RESET, A2 => n2387, ZN => n2470);
   U1837 : OAI21_X1 port map( B1 => n3582, B2 => n2473, A => n2474, ZN => n1731
                           );
   U1838 : MUX2_X1 port map( A => n3515, B => n2475, S => n2476, Z => 
                           n1730_port);
   U1839 : MUX2_X1 port map( A => n3514, B => n2477, S => n2476, Z => 
                           n1729_port);
   U1840 : MUX2_X1 port map( A => n3513, B => n2478, S => n2476, Z => 
                           n1728_port);
   U1841 : MUX2_X1 port map( A => n3512, B => n2479, S => n2476, Z => 
                           n1727_port);
   U1842 : MUX2_X1 port map( A => n3511, B => n2480, S => n2476, Z => 
                           n1726_port);
   U1843 : MUX2_X1 port map( A => n3510, B => n2481, S => n2476, Z => 
                           n1725_port);
   U1844 : MUX2_X1 port map( A => n3509, B => n2482, S => n2476, Z => n1724);
   U1845 : MUX2_X1 port map( A => n3508, B => n2483, S => n2476, Z => n1723);
   U1846 : OAI221_X1 port map( B1 => n2484, B2 => n2485, C1 => n2486, C2 => 
                           n2487, A => n2374, ZN => n2476);
   U1847 : MUX2_X1 port map( A => n3507, B => n2475, S => n2488, Z => n1722);
   U1848 : MUX2_X1 port map( A => n3506, B => n2477, S => n2488, Z => n1721);
   U1849 : MUX2_X1 port map( A => n3505, B => n2478, S => n2488, Z => n1720);
   U1850 : MUX2_X1 port map( A => n3504, B => n2479, S => n2488, Z => n1719);
   U1851 : MUX2_X1 port map( A => n3503, B => n2480, S => n2488, Z => n1718);
   U1852 : MUX2_X1 port map( A => n3502, B => n2481, S => n2488, Z => n1717);
   U1853 : MUX2_X1 port map( A => n3501, B => n2482, S => n2488, Z => n1716);
   U1854 : MUX2_X1 port map( A => n3500, B => n2483, S => n2488, Z => n1715);
   U1855 : OAI221_X1 port map( B1 => n2485, B2 => n2489, C1 => n2486, C2 => 
                           n2490, A => n2374, ZN => n2488);
   U1856 : MUX2_X1 port map( A => n3499, B => n2475, S => n2491, Z => n1714);
   U1857 : MUX2_X1 port map( A => n3498, B => n2477, S => n2491, Z => n1713);
   U1858 : MUX2_X1 port map( A => n3497, B => n2478, S => n2491, Z => n1712);
   U1859 : MUX2_X1 port map( A => n3496, B => n2479, S => n2491, Z => n1711);
   U1860 : MUX2_X1 port map( A => n3495, B => n2480, S => n2491, Z => n1710);
   U1861 : MUX2_X1 port map( A => n3494, B => n2481, S => n2491, Z => n1709);
   U1862 : MUX2_X1 port map( A => n3493, B => n2482, S => n2491, Z => n1708);
   U1863 : MUX2_X1 port map( A => n3492, B => n2483, S => n2491, Z => n1707);
   U1864 : OAI221_X1 port map( B1 => n2485, B2 => n2492, C1 => n2472, C2 => 
                           n2493, A => n2374, ZN => n2491);
   U1865 : MUX2_X1 port map( A => n3491, B => n2475, S => n2494, Z => n1706);
   U1866 : MUX2_X1 port map( A => n3490, B => n2477, S => n2494, Z => n1705);
   U1867 : MUX2_X1 port map( A => n3489, B => n2478, S => n2494, Z => n1704);
   U1868 : MUX2_X1 port map( A => n3488, B => n2479, S => n2494, Z => n1703);
   U1869 : MUX2_X1 port map( A => n3487, B => n2480, S => n2494, Z => n1702);
   U1870 : MUX2_X1 port map( A => n3486, B => n2481, S => n2494, Z => n1701);
   U1871 : MUX2_X1 port map( A => n3485, B => n2482, S => n2494, Z => n1700);
   U1872 : MUX2_X1 port map( A => n3484, B => n2483, S => n2494, Z => n1699);
   U1873 : OAI221_X1 port map( B1 => n2485, B2 => n2495, C1 => n2472, C2 => 
                           n2496, A => n2374, ZN => n2494);
   U1874 : MUX2_X1 port map( A => n3483, B => n2475, S => n2497, Z => n1698);
   U1875 : MUX2_X1 port map( A => n3482, B => n2477, S => n2497, Z => n1697);
   U1876 : MUX2_X1 port map( A => n3481, B => n2478, S => n2497, Z => n1696);
   U1877 : MUX2_X1 port map( A => n3480, B => n2479, S => n2497, Z => n1695);
   U1878 : MUX2_X1 port map( A => n3479, B => n2480, S => n2497, Z => n1694);
   U1879 : MUX2_X1 port map( A => n3478, B => n2481, S => n2497, Z => n1693);
   U1880 : MUX2_X1 port map( A => n3477, B => n2482, S => n2497, Z => n1692);
   U1881 : MUX2_X1 port map( A => n3476, B => n2483, S => n2497, Z => n1691);
   U1882 : OAI221_X1 port map( B1 => n2498, B2 => n2499, C1 => n2484, C2 => 
                           n2500, A => n2374, ZN => n2497);
   U1883 : MUX2_X1 port map( A => n3475, B => n2475, S => n2501, Z => n1690);
   U1884 : MUX2_X1 port map( A => n3474, B => n2477, S => n2501, Z => n1689);
   U1885 : MUX2_X1 port map( A => n3473, B => n2478, S => n2501, Z => n1688);
   U1886 : MUX2_X1 port map( A => n3472, B => n2479, S => n2501, Z => n1687);
   U1887 : MUX2_X1 port map( A => n3471, B => n2480, S => n2501, Z => n1686);
   U1888 : MUX2_X1 port map( A => n3470, B => n2481, S => n2501, Z => n1685);
   U1889 : MUX2_X1 port map( A => n3469, B => n2482, S => n2501, Z => n1684);
   U1890 : MUX2_X1 port map( A => n3468, B => n2483, S => n2501, Z => n1683);
   U1891 : OAI221_X1 port map( B1 => n2499, B2 => n2502, C1 => n2489, C2 => 
                           n2500, A => n2374, ZN => n2501);
   U1892 : MUX2_X1 port map( A => n3467, B => n2475, S => n2503, Z => n1682);
   U1893 : MUX2_X1 port map( A => n3466, B => n2477, S => n2503, Z => n1681);
   U1894 : MUX2_X1 port map( A => n3465, B => n2478, S => n2503, Z => n1680);
   U1895 : MUX2_X1 port map( A => n3464, B => n2479, S => n2503, Z => n1679);
   U1896 : MUX2_X1 port map( A => n3463, B => n2480, S => n2503, Z => n1678);
   U1897 : MUX2_X1 port map( A => n3462, B => n2481, S => n2503, Z => n1677);
   U1898 : MUX2_X1 port map( A => n3461, B => n2482, S => n2503, Z => n1676);
   U1899 : MUX2_X1 port map( A => n3460, B => n2483, S => n2503, Z => n1675);
   U1900 : OAI221_X1 port map( B1 => n2492, B2 => n2500, C1 => n2472, C2 => 
                           n2504, A => n2374, ZN => n2503);
   U1901 : MUX2_X1 port map( A => n3459, B => n2475, S => n2505, Z => n1674);
   U1902 : MUX2_X1 port map( A => n3458, B => n2477, S => n2505, Z => n1673);
   U1903 : MUX2_X1 port map( A => n3457, B => n2478, S => n2505, Z => n1672);
   U1904 : MUX2_X1 port map( A => n3456, B => n2479, S => n2505, Z => n1671);
   U1905 : MUX2_X1 port map( A => n3455, B => n2480, S => n2505, Z => n1670);
   U1906 : MUX2_X1 port map( A => n3454, B => n2481, S => n2505, Z => n1669);
   U1907 : MUX2_X1 port map( A => n3453, B => n2482, S => n2505, Z => n1668);
   U1908 : MUX2_X1 port map( A => n3452, B => n2483, S => n2505, Z => n1667);
   U1909 : OAI221_X1 port map( B1 => n2495, B2 => n2500, C1 => n2472, C2 => 
                           n2506, A => n2374, ZN => n2505);
   U1910 : MUX2_X1 port map( A => n3451, B => n2475, S => n2507, Z => n1666);
   U1911 : MUX2_X1 port map( A => n3450, B => n2477, S => n2507, Z => n1665);
   U1912 : MUX2_X1 port map( A => n3449, B => n2478, S => n2507, Z => n1664);
   U1913 : MUX2_X1 port map( A => n3448, B => n2479, S => n2507, Z => n1663);
   U1914 : MUX2_X1 port map( A => n3447, B => n2480, S => n2507, Z => n1662);
   U1915 : MUX2_X1 port map( A => n3446, B => n2481, S => n2507, Z => n1661);
   U1916 : MUX2_X1 port map( A => n3445, B => n2482, S => n2507, Z => n1660);
   U1917 : MUX2_X1 port map( A => n3444, B => n2483, S => n2507, Z => n1659);
   U1918 : OAI221_X1 port map( B1 => n2498, B2 => n2508, C1 => n2484, C2 => 
                           n2509, A => n2374, ZN => n2507);
   U1919 : MUX2_X1 port map( A => n3443, B => n2475, S => n2510, Z => n1658);
   U1920 : MUX2_X1 port map( A => n3442, B => n2477, S => n2510, Z => n1657);
   U1921 : MUX2_X1 port map( A => n3441, B => n2478, S => n2510, Z => n1656);
   U1922 : MUX2_X1 port map( A => n3440, B => n2479, S => n2510, Z => n1655);
   U1923 : MUX2_X1 port map( A => n3439, B => n2480, S => n2510, Z => n1654);
   U1924 : MUX2_X1 port map( A => n3438, B => n2481, S => n2510, Z => n1653);
   U1925 : MUX2_X1 port map( A => n3437, B => n2482, S => n2510, Z => n1652);
   U1926 : MUX2_X1 port map( A => n3436, B => n2483, S => n2510, Z => n1651);
   U1927 : OAI221_X1 port map( B1 => n2502, B2 => n2508, C1 => n2489, C2 => 
                           n2509, A => n2374, ZN => n2510);
   U1928 : MUX2_X1 port map( A => n3435, B => n2475, S => n2511, Z => n1650);
   U1929 : MUX2_X1 port map( A => n3434, B => n2477, S => n2511, Z => n1649);
   U1930 : MUX2_X1 port map( A => n3433, B => n2478, S => n2511, Z => n1648);
   U1931 : MUX2_X1 port map( A => n3432, B => n2479, S => n2511, Z => n1647);
   U1932 : MUX2_X1 port map( A => n3431, B => n2480, S => n2511, Z => n1646);
   U1933 : MUX2_X1 port map( A => n3430, B => n2481, S => n2511, Z => n1645);
   U1934 : MUX2_X1 port map( A => n3429, B => n2482, S => n2511, Z => n1644);
   U1935 : MUX2_X1 port map( A => n3428, B => n2483, S => n2511, Z => n1643);
   U1936 : OAI221_X1 port map( B1 => n2492, B2 => n2509, C1 => n2472, C2 => 
                           n2512, A => n2374, ZN => n2511);
   U1937 : MUX2_X1 port map( A => n3427, B => n2475, S => n2513, Z => n1642);
   U1938 : MUX2_X1 port map( A => n3426, B => n2477, S => n2513, Z => n1641);
   U1939 : MUX2_X1 port map( A => n3425, B => n2478, S => n2513, Z => n1640);
   U1940 : MUX2_X1 port map( A => n3424, B => n2479, S => n2513, Z => n1639);
   U1941 : MUX2_X1 port map( A => n3423, B => n2480, S => n2513, Z => n1638);
   U1942 : MUX2_X1 port map( A => n3422, B => n2481, S => n2513, Z => n1637);
   U1943 : MUX2_X1 port map( A => n3421, B => n2482, S => n2513, Z => n1636);
   U1944 : MUX2_X1 port map( A => n3420, B => n2483, S => n2513, Z => n1635);
   U1945 : OAI221_X1 port map( B1 => n2495, B2 => n2509, C1 => n2472, C2 => 
                           n2514, A => n2374, ZN => n2513);
   U1946 : MUX2_X1 port map( A => n3419, B => n2475, S => n2515, Z => n1634);
   U1947 : MUX2_X1 port map( A => n3418, B => n2477, S => n2515, Z => n1633);
   U1948 : MUX2_X1 port map( A => n3417, B => n2478, S => n2515, Z => n1632);
   U1949 : MUX2_X1 port map( A => n3416, B => n2479, S => n2515, Z => n1631);
   U1950 : MUX2_X1 port map( A => n3415, B => n2480, S => n2515, Z => n1630);
   U1951 : MUX2_X1 port map( A => n3414, B => n2481, S => n2515, Z => n1629);
   U1952 : MUX2_X1 port map( A => n3413, B => n2482, S => n2515, Z => n1628);
   U1953 : MUX2_X1 port map( A => n3412, B => n2483, S => n2515, Z => n1627);
   U1954 : OAI221_X1 port map( B1 => n2498, B2 => n2516, C1 => n2484, C2 => 
                           n2517, A => n2374, ZN => n2515);
   U1955 : NAND3_X1 port map( A1 => n2420, A2 => n2421, A3 => n2518, ZN => 
                           n2484);
   U1956 : NAND2_X1 port map( A1 => n2519, A2 => n2080, ZN => n2498);
   U1957 : MUX2_X1 port map( A => n3411, B => n2475, S => n2520, Z => n1626);
   U1958 : MUX2_X1 port map( A => n3410, B => n2477, S => n2520, Z => n1625);
   U1959 : MUX2_X1 port map( A => n3409, B => n2478, S => n2520, Z => n1624);
   U1960 : MUX2_X1 port map( A => n3408, B => n2479, S => n2520, Z => n1623);
   U1961 : MUX2_X1 port map( A => n3407, B => n2480, S => n2520, Z => n1622);
   U1962 : MUX2_X1 port map( A => n3406, B => n2481, S => n2520, Z => n1621);
   U1963 : MUX2_X1 port map( A => n3405, B => n2482, S => n2520, Z => n1620);
   U1964 : MUX2_X1 port map( A => n3404, B => n2483, S => n2520, Z => n1619);
   U1965 : OAI221_X1 port map( B1 => n2502, B2 => n2516, C1 => n2489, C2 => 
                           n2517, A => n2374, ZN => n2520);
   U1966 : NAND3_X1 port map( A1 => N302, A2 => n2421, A3 => n2518, ZN => n2489
                           );
   U1967 : NAND2_X1 port map( A1 => n2521, A2 => n2080, ZN => n2502);
   U1968 : MUX2_X1 port map( A => n3403, B => n2475, S => n2522, Z => n1618);
   U1969 : MUX2_X1 port map( A => n3402, B => n2477, S => n2522, Z => n1617);
   U1970 : MUX2_X1 port map( A => n3401, B => n2478, S => n2522, Z => n1616);
   U1971 : MUX2_X1 port map( A => n3400, B => n2479, S => n2522, Z => n1615);
   U1972 : MUX2_X1 port map( A => n3399, B => n2480, S => n2522, Z => n1614);
   U1973 : MUX2_X1 port map( A => n3398, B => n2481, S => n2522, Z => n1613);
   U1974 : MUX2_X1 port map( A => n3397, B => n2482, S => n2522, Z => n1612);
   U1975 : MUX2_X1 port map( A => n3396, B => n2483, S => n2522, Z => n1611);
   U1976 : OAI221_X1 port map( B1 => n2492, B2 => n2517, C1 => n2472, C2 => 
                           n2523, A => n2374, ZN => n2522);
   U1977 : NAND3_X1 port map( A1 => N303, A2 => n2420, A3 => n2518, ZN => n2492
                           );
   U1978 : MUX2_X1 port map( A => n3395, B => n2475, S => n2524, Z => n1610);
   U1979 : MUX2_X1 port map( A => n3394, B => n2477, S => n2524, Z => n1609);
   U1980 : MUX2_X1 port map( A => n3393, B => n2478, S => n2524, Z => n1608);
   U1981 : MUX2_X1 port map( A => n3392, B => n2479, S => n2524, Z => n1607);
   U1982 : MUX2_X1 port map( A => n3391, B => n2480, S => n2524, Z => n1606);
   U1983 : MUX2_X1 port map( A => n3390, B => n2481, S => n2524, Z => n1605);
   U1984 : MUX2_X1 port map( A => n3389, B => n2482, S => n2524, Z => n1604);
   U1985 : MUX2_X1 port map( A => n3388, B => n2483, S => n2524, Z => n1603);
   U1986 : OAI221_X1 port map( B1 => n2495, B2 => n2517, C1 => n2472, C2 => 
                           n2525, A => n2374, ZN => n2524);
   U1987 : NAND3_X1 port map( A1 => N303, A2 => N302, A3 => n2518, ZN => n2495)
                           ;
   U1988 : AND4_X1 port map( A1 => WR, A2 => n2432, A3 => n2526, A4 => n2527, 
                           ZN => n2518);
   U1989 : INV_X1 port map( A => N312, ZN => n2527);
   U1990 : MUX2_X1 port map( A => n3387, B => n2475, S => n2528, Z => n1602);
   U1991 : MUX2_X1 port map( A => n3386, B => n2477, S => n2528, Z => n1601);
   U1992 : MUX2_X1 port map( A => n3385, B => n2478, S => n2528, Z => n1600);
   U1993 : MUX2_X1 port map( A => n3384, B => n2479, S => n2528, Z => n1599);
   U1994 : MUX2_X1 port map( A => n3383, B => n2480, S => n2528, Z => n1598);
   U1995 : MUX2_X1 port map( A => n3382, B => n2481, S => n2528, Z => n1597);
   U1996 : MUX2_X1 port map( A => n3381, B => n2482, S => n2528, Z => n1596);
   U1997 : MUX2_X1 port map( A => n3380, B => n2483, S => n2528, Z => n1595);
   U1998 : OAI221_X1 port map( B1 => n2485, B2 => n2529, C1 => n2487, C2 => 
                           n2530, A => n2374, ZN => n2528);
   U1999 : INV_X1 port map( A => n2519, ZN => n2487);
   U2000 : MUX2_X1 port map( A => n3379, B => n2475, S => n2531, Z => n1594);
   U2001 : MUX2_X1 port map( A => n3378, B => n2477, S => n2531, Z => n1593);
   U2002 : MUX2_X1 port map( A => n3377, B => n2478, S => n2531, Z => n1592);
   U2003 : MUX2_X1 port map( A => n3376, B => n2479, S => n2531, Z => n1591);
   U2004 : MUX2_X1 port map( A => n3375, B => n2480, S => n2531, Z => n1590);
   U2005 : MUX2_X1 port map( A => n3374, B => n2481, S => n2531, Z => n1589);
   U2006 : MUX2_X1 port map( A => n3373, B => n2482, S => n2531, Z => n1588);
   U2007 : MUX2_X1 port map( A => n3372, B => n2483, S => n2531, Z => n1587);
   U2008 : OAI221_X1 port map( B1 => n2485, B2 => n2532, C1 => n2490, C2 => 
                           n2530, A => n2374, ZN => n2531);
   U2009 : INV_X1 port map( A => n2521, ZN => n2490);
   U2010 : MUX2_X1 port map( A => n3371, B => n2475, S => n2533, Z => n1586);
   U2011 : MUX2_X1 port map( A => n3370, B => n2477, S => n2533, Z => n1585);
   U2012 : MUX2_X1 port map( A => n3369, B => n2478, S => n2533, Z => n1584);
   U2013 : MUX2_X1 port map( A => n3368, B => n2479, S => n2533, Z => n1583);
   U2014 : MUX2_X1 port map( A => n3367, B => n2480, S => n2533, Z => n1582);
   U2015 : MUX2_X1 port map( A => n3366, B => n2481, S => n2533, Z => n1581);
   U2016 : MUX2_X1 port map( A => n3365, B => n2482, S => n2533, Z => n1580);
   U2017 : MUX2_X1 port map( A => n3364, B => n2483, S => n2533, Z => n1579);
   U2018 : OAI221_X1 port map( B1 => n2485, B2 => n2534, C1 => n2472, C2 => 
                           n2535, A => n2374, ZN => n2533);
   U2019 : MUX2_X1 port map( A => n3363, B => n2475, S => n2536, Z => n1578);
   U2020 : MUX2_X1 port map( A => n3362, B => n2477, S => n2536, Z => n1577);
   U2021 : MUX2_X1 port map( A => n3361, B => n2478, S => n2536, Z => n1576);
   U2022 : MUX2_X1 port map( A => n3360, B => n2479, S => n2536, Z => n1575);
   U2023 : MUX2_X1 port map( A => n3359, B => n2480, S => n2536, Z => n1574);
   U2024 : MUX2_X1 port map( A => n3358, B => n2481, S => n2536, Z => n1573);
   U2025 : MUX2_X1 port map( A => n3357, B => n2482, S => n2536, Z => n1572);
   U2026 : MUX2_X1 port map( A => n3356, B => n2483, S => n2536, Z => n1571);
   U2027 : OAI221_X1 port map( B1 => n2485, B2 => n2537, C1 => n2472, C2 => 
                           n2538, A => n2374, ZN => n2536);
   U2028 : NAND2_X1 port map( A1 => n2539, A2 => n2540, ZN => n2485);
   U2029 : MUX2_X1 port map( A => n3355, B => n2475, S => n2541, Z => n1570);
   U2030 : MUX2_X1 port map( A => n3354, B => n2477, S => n2541, Z => n1569);
   U2031 : MUX2_X1 port map( A => n3353, B => n2478, S => n2541, Z => n1568);
   U2032 : MUX2_X1 port map( A => n3352, B => n2479, S => n2541, Z => n1567);
   U2033 : MUX2_X1 port map( A => n3351, B => n2480, S => n2541, Z => n1566);
   U2034 : MUX2_X1 port map( A => n3350, B => n2481, S => n2541, Z => n1565);
   U2035 : MUX2_X1 port map( A => n3349, B => n2482, S => n2541, Z => n1564);
   U2036 : MUX2_X1 port map( A => n3348, B => n2483, S => n2541, Z => n1563);
   U2037 : OAI221_X1 port map( B1 => n2499, B2 => n2542, C1 => n2500, C2 => 
                           n2529, A => n2374, ZN => n2541);
   U2038 : MUX2_X1 port map( A => n3347, B => n2475, S => n2543, Z => n1562);
   U2039 : MUX2_X1 port map( A => n3346, B => n2477, S => n2543, Z => n1561);
   U2040 : MUX2_X1 port map( A => n3345, B => n2478, S => n2543, Z => n1560);
   U2041 : MUX2_X1 port map( A => n3344, B => n2479, S => n2543, Z => n1559);
   U2042 : MUX2_X1 port map( A => n3343, B => n2480, S => n2543, Z => n1558);
   U2043 : MUX2_X1 port map( A => n3342, B => n2481, S => n2543, Z => n1557);
   U2044 : MUX2_X1 port map( A => n3341, B => n2482, S => n2543, Z => n1556);
   U2045 : MUX2_X1 port map( A => n3340, B => n2483, S => n2543, Z => n1555);
   U2046 : OAI221_X1 port map( B1 => n2499, B2 => n2544, C1 => n2500, C2 => 
                           n2532, A => n2374, ZN => n2543);
   U2047 : MUX2_X1 port map( A => n3339, B => n2475, S => n2545, Z => n1554);
   U2048 : MUX2_X1 port map( A => n3338, B => n2477, S => n2545, Z => n1553);
   U2049 : MUX2_X1 port map( A => n3337, B => n2478, S => n2545, Z => n1552);
   U2050 : MUX2_X1 port map( A => n3336, B => n2479, S => n2545, Z => n1551);
   U2051 : MUX2_X1 port map( A => n3335, B => n2480, S => n2545, Z => n1550);
   U2052 : MUX2_X1 port map( A => n3334, B => n2481, S => n2545, Z => n1549);
   U2053 : MUX2_X1 port map( A => n3333, B => n2482, S => n2545, Z => n1548);
   U2054 : MUX2_X1 port map( A => n3332, B => n2483, S => n2545, Z => n1547);
   U2055 : OAI221_X1 port map( B1 => n2500, B2 => n2534, C1 => n2472, C2 => 
                           n2546, A => n2374, ZN => n2545);
   U2056 : MUX2_X1 port map( A => n3331, B => n2475, S => n2547, Z => n1546);
   U2057 : MUX2_X1 port map( A => n3330, B => n2477, S => n2547, Z => n1545);
   U2058 : MUX2_X1 port map( A => n3329, B => n2478, S => n2547, Z => n1544);
   U2059 : MUX2_X1 port map( A => n3328, B => n2479, S => n2547, Z => n1543);
   U2060 : MUX2_X1 port map( A => n3327, B => n2480, S => n2547, Z => n1542);
   U2061 : MUX2_X1 port map( A => n3326, B => n2481, S => n2547, Z => n1541);
   U2062 : MUX2_X1 port map( A => n3325, B => n2482, S => n2547, Z => n1540);
   U2063 : MUX2_X1 port map( A => n3324, B => n2483, S => n2547, Z => n1539);
   U2064 : OAI221_X1 port map( B1 => n2500, B2 => n2537, C1 => n2472, C2 => 
                           n2548, A => n2374, ZN => n2547);
   U2065 : NAND2_X1 port map( A1 => N310, A2 => n2539, ZN => n2500);
   U2066 : INV_X1 port map( A => N311, ZN => n2539);
   U2067 : MUX2_X1 port map( A => n3323, B => n2475, S => n2549, Z => n1538);
   U2068 : MUX2_X1 port map( A => n3322, B => n2477, S => n2549, Z => n1537);
   U2069 : MUX2_X1 port map( A => n3321, B => n2478, S => n2549, Z => n1536);
   U2070 : MUX2_X1 port map( A => n3320, B => n2479, S => n2549, Z => n1535);
   U2071 : MUX2_X1 port map( A => n3319, B => n2480, S => n2549, Z => n1534);
   U2072 : MUX2_X1 port map( A => n3318, B => n2481, S => n2549, Z => n1533);
   U2073 : MUX2_X1 port map( A => n3317, B => n2482, S => n2549, Z => n1532);
   U2074 : MUX2_X1 port map( A => n3316, B => n2483, S => n2549, Z => n1531);
   U2075 : OAI221_X1 port map( B1 => n2508, B2 => n2542, C1 => n2509, C2 => 
                           n2529, A => n2374, ZN => n2549);
   U2076 : MUX2_X1 port map( A => n3315, B => n2475, S => n2550, Z => n1530);
   U2077 : MUX2_X1 port map( A => n3314, B => n2477, S => n2550, Z => n1529);
   U2078 : MUX2_X1 port map( A => n3313, B => n2478, S => n2550, Z => n1528);
   U2079 : MUX2_X1 port map( A => n3312, B => n2479, S => n2550, Z => n1527);
   U2080 : MUX2_X1 port map( A => n3311, B => n2480, S => n2550, Z => n1526);
   U2081 : MUX2_X1 port map( A => n3310, B => n2481, S => n2550, Z => n1525);
   U2082 : MUX2_X1 port map( A => n3309, B => n2482, S => n2550, Z => n1524);
   U2083 : MUX2_X1 port map( A => n3308, B => n2483, S => n2550, Z => n1523);
   U2084 : OAI221_X1 port map( B1 => n2508, B2 => n2544, C1 => n2509, C2 => 
                           n2532, A => n2374, ZN => n2550);
   U2085 : MUX2_X1 port map( A => n3307, B => n2475, S => n2551, Z => n1522);
   U2086 : MUX2_X1 port map( A => n3306, B => n2477, S => n2551, Z => n1521);
   U2087 : MUX2_X1 port map( A => n3305, B => n2478, S => n2551, Z => n1520);
   U2088 : MUX2_X1 port map( A => n3304, B => n2479, S => n2551, Z => n1519);
   U2089 : MUX2_X1 port map( A => n3303, B => n2480, S => n2551, Z => n1518);
   U2090 : MUX2_X1 port map( A => n3302, B => n2481, S => n2551, Z => n1517);
   U2091 : MUX2_X1 port map( A => n3301, B => n2482, S => n2551, Z => n1516);
   U2092 : MUX2_X1 port map( A => n3300, B => n2483, S => n2551, Z => n1515);
   U2093 : OAI221_X1 port map( B1 => n2509, B2 => n2534, C1 => n2472, C2 => 
                           n2552, A => n2374, ZN => n2551);
   U2094 : MUX2_X1 port map( A => n3299, B => n2475, S => n2553, Z => n1514);
   U2095 : MUX2_X1 port map( A => n3298, B => n2477, S => n2553, Z => n1513);
   U2096 : MUX2_X1 port map( A => n3297, B => n2478, S => n2553, Z => n1512);
   U2097 : MUX2_X1 port map( A => n3296, B => n2479, S => n2553, Z => n1511);
   U2098 : MUX2_X1 port map( A => n3295, B => n2480, S => n2553, Z => n1510);
   U2099 : MUX2_X1 port map( A => n3294, B => n2481, S => n2553, Z => n1509);
   U2100 : MUX2_X1 port map( A => n3293, B => n2482, S => n2553, Z => n1508);
   U2101 : MUX2_X1 port map( A => n3292, B => n2483, S => n2553, Z => n1507);
   U2102 : OAI221_X1 port map( B1 => n2509, B2 => n2537, C1 => n2472, C2 => 
                           n2554, A => n2374, ZN => n2553);
   U2103 : NAND2_X1 port map( A1 => N311, A2 => n2540, ZN => n2509);
   U2104 : INV_X1 port map( A => N310, ZN => n2540);
   U2105 : MUX2_X1 port map( A => n3291, B => n2475, S => n2555, Z => n1506);
   U2106 : MUX2_X1 port map( A => n3290, B => n2477, S => n2555, Z => n1505);
   U2107 : MUX2_X1 port map( A => n3289, B => n2478, S => n2555, Z => n1504);
   U2108 : MUX2_X1 port map( A => n3288, B => n2479, S => n2555, Z => n1503);
   U2109 : MUX2_X1 port map( A => n3287, B => n2480, S => n2555, Z => n1502);
   U2110 : MUX2_X1 port map( A => n3286, B => n2481, S => n2555, Z => n1501);
   U2111 : MUX2_X1 port map( A => n3285, B => n2482, S => n2555, Z => n1500);
   U2112 : MUX2_X1 port map( A => n3284, B => n2483, S => n2555, Z => n1499);
   U2113 : OAI221_X1 port map( B1 => n2516, B2 => n2542, C1 => n2517, C2 => 
                           n2529, A => n2374, ZN => n2555);
   U2114 : NAND3_X1 port map( A1 => n2420, A2 => n2421, A3 => n2556, ZN => 
                           n2529);
   U2115 : NAND2_X1 port map( A1 => n2519, A2 => n3585, ZN => n2542);
   U2116 : NOR2_X1 port map( A1 => n2472, A2 => n2557, ZN => n2519);
   U2117 : MUX2_X1 port map( A => n3283, B => n2475, S => n2558, Z => n1498);
   U2118 : MUX2_X1 port map( A => n3282, B => n2477, S => n2558, Z => n1497);
   U2119 : MUX2_X1 port map( A => n3281, B => n2478, S => n2558, Z => n1496);
   U2120 : MUX2_X1 port map( A => n3280, B => n2479, S => n2558, Z => n1495);
   U2121 : MUX2_X1 port map( A => n3279, B => n2480, S => n2558, Z => n1494);
   U2122 : MUX2_X1 port map( A => n3278, B => n2481, S => n2558, Z => n1493);
   U2123 : MUX2_X1 port map( A => n3277, B => n2482, S => n2558, Z => n1492);
   U2124 : MUX2_X1 port map( A => n3276, B => n2483, S => n2558, Z => n1491);
   U2125 : OAI221_X1 port map( B1 => n2516, B2 => n2544, C1 => n2517, C2 => 
                           n2532, A => n2374, ZN => n2558);
   U2126 : NAND3_X1 port map( A1 => N302, A2 => n2421, A3 => n2556, ZN => n2532
                           );
   U2127 : INV_X1 port map( A => N303, ZN => n2421);
   U2128 : NAND2_X1 port map( A1 => n2521, A2 => n3585, ZN => n2544);
   U2129 : NOR3_X1 port map( A1 => n2188, A2 => n3588, A3 => n2472, ZN => n2521
                           );
   U2130 : MUX2_X1 port map( A => n2190, B => n2475, S => n2559, Z => n1490);
   U2131 : MUX2_X1 port map( A => n2192, B => n2477, S => n2559, Z => n1489);
   U2132 : MUX2_X1 port map( A => n2194, B => n2478, S => n2559, Z => n1488);
   U2133 : MUX2_X1 port map( A => n2196, B => n2479, S => n2559, Z => n1487);
   U2134 : MUX2_X1 port map( A => n2197, B => n2480, S => n2559, Z => n1486);
   U2135 : MUX2_X1 port map( A => n2195, B => n2481, S => n2559, Z => n1485);
   U2136 : MUX2_X1 port map( A => n2193, B => n2482, S => n2559, Z => n1484);
   U2137 : MUX2_X1 port map( A => n2191, B => n2483, S => n2559, Z => n1483);
   U2138 : OAI221_X1 port map( B1 => n2517, B2 => n2534, C1 => n2472, C2 => 
                           n2560, A => n2374, ZN => n2559);
   U2139 : NAND3_X1 port map( A1 => N303, A2 => n2420, A3 => n2556, ZN => n2534
                           );
   U2140 : INV_X1 port map( A => N302, ZN => n2420);
   U2141 : MUX2_X1 port map( A => n2083, B => n2475, S => n2561, Z => n1482);
   U2142 : AND2_X1 port map( A1 => n2562, A2 => n2374, ZN => n2475);
   U2143 : MUX2_X1 port map( A => DATA_FROM_MEM(7), B => DATAIN(7), S => n2389,
                           Z => n2562);
   U2144 : MUX2_X1 port map( A => n2085, B => n2477, S => n2561, Z => n1481);
   U2145 : AND2_X1 port map( A1 => n2563, A2 => n2374, ZN => n2477);
   U2146 : MUX2_X1 port map( A => DATA_FROM_MEM(5), B => DATAIN(5), S => n2389,
                           Z => n2563);
   U2147 : MUX2_X1 port map( A => n2087, B => n2478, S => n2561, Z => n1480);
   U2148 : AND2_X1 port map( A1 => n2564, A2 => n2374, ZN => n2478);
   U2149 : MUX2_X1 port map( A => DATA_FROM_MEM(3), B => DATAIN(3), S => n2389,
                           Z => n2564);
   U2150 : MUX2_X1 port map( A => n2089, B => n2479, S => n2561, Z => n1479);
   U2151 : AND2_X1 port map( A1 => n2565, A2 => n2374, ZN => n2479);
   U2152 : MUX2_X1 port map( A => DATA_FROM_MEM(1), B => DATAIN(1), S => n2389,
                           Z => n2565);
   U2153 : MUX2_X1 port map( A => n2090, B => n2480, S => n2561, Z => n1478);
   U2154 : AND2_X1 port map( A1 => n2566, A2 => n2374, ZN => n2480);
   U2155 : MUX2_X1 port map( A => DATA_FROM_MEM(0), B => DATAIN(0), S => n2389,
                           Z => n2566);
   U2156 : MUX2_X1 port map( A => n2088, B => n2481, S => n2561, Z => n1477);
   U2157 : AND2_X1 port map( A1 => n2567, A2 => n2374, ZN => n2481);
   U2158 : MUX2_X1 port map( A => DATA_FROM_MEM(2), B => DATAIN(2), S => n2389,
                           Z => n2567);
   U2159 : MUX2_X1 port map( A => n2086, B => n2482, S => n2561, Z => n1476);
   U2160 : AND2_X1 port map( A1 => n2568, A2 => n2374, ZN => n2482);
   U2161 : MUX2_X1 port map( A => DATA_FROM_MEM(4), B => DATAIN(4), S => n2389,
                           Z => n2568);
   U2162 : MUX2_X1 port map( A => n2084, B => n2483, S => n2561, Z => n1475);
   U2163 : OAI221_X1 port map( B1 => n2472, B2 => n2569, C1 => n2517, C2 => 
                           n2537, A => n2374, ZN => n2561);
   U2164 : NAND3_X1 port map( A1 => N303, A2 => N302, A3 => n2556, ZN => n2537)
                           ;
   U2165 : AND4_X1 port map( A1 => N312, A2 => WR, A3 => n2432, A4 => n2526, ZN
                           => n2556);
   U2166 : NAND2_X1 port map( A1 => N311, A2 => N310, ZN => n2517);
   U2167 : NAND2_X1 port map( A1 => n2570, A2 => ENABLE, ZN => n2472);
   U2168 : AND2_X1 port map( A1 => n2571, A2 => n2374, ZN => n2483);
   U2169 : MUX2_X1 port map( A => DATA_FROM_MEM(6), B => DATAIN(6), S => n2389,
                           Z => n2571);
   U2170 : OAI211_X1 port map( C1 => n2572, C2 => n2352, A => n2573, B => n2574
                           , ZN => n1474);
   U2171 : AOI221_X1 port map( B1 => n2575, B2 => n3531, C1 => n2576, C2 => 
                           n2231, A => n2577, ZN => n2574);
   U2172 : AOI21_X1 port map( B1 => n2578, B2 => n2579, A => n2580, ZN => n2577
                           );
   U2173 : NOR4_X1 port map( A1 => n2581, A2 => n2582, A3 => n2583, A4 => n2584
                           , ZN => n2579);
   U2174 : OAI221_X1 port map( B1 => n2131, B2 => n2585, C1 => n2248, C2 => 
                           n2586, A => n2587, ZN => n2584);
   U2175 : AOI22_X1 port map( A1 => n2588, A2 => n3411, B1 => n2589, B2 => 
                           n3419, ZN => n2587);
   U2176 : OAI221_X1 port map( B1 => n2132, B2 => n2590, C1 => n2256, C2 => 
                           n2591, A => n2592, ZN => n2583);
   U2177 : AOI22_X1 port map( A1 => n2593, A2 => n3475, B1 => n2594, B2 => 
                           n3483, ZN => n2592);
   U2178 : OAI221_X1 port map( B1 => n2107, B2 => n2595, C1 => n2198, C2 => 
                           n2596, A => n2597, ZN => n2582);
   U2179 : AOI22_X1 port map( A1 => n2598, A2 => n2083, B1 => n2599, B2 => 
                           n2190, ZN => n2597);
   U2180 : OAI221_X1 port map( B1 => n2108, B2 => n2600, C1 => n2199, C2 => 
                           n2601, A => n2602, ZN => n2581);
   U2181 : AOI22_X1 port map( A1 => n2603, A2 => n3379, B1 => n2604, B2 => 
                           n3387, ZN => n2602);
   U2182 : NOR4_X1 port map( A1 => n2605, A2 => n2606, A3 => n2607, A4 => n2608
                           , ZN => n2578);
   U2183 : OAI221_X1 port map( B1 => n2123, B2 => n2609, C1 => n2272, C2 => 
                           n2610, A => n2611, ZN => n2608);
   U2184 : AOI22_X1 port map( A1 => n2612, A2 => n3435, B1 => n2613, B2 => 
                           n3427, ZN => n2611);
   U2185 : OAI221_X1 port map( B1 => n2147, B2 => n2614, C1 => n2264, C2 => 
                           n2615, A => n2616, ZN => n2607);
   U2186 : AOI22_X1 port map( A1 => n2617, A2 => n3499, B1 => n2618, B2 => 
                           n3491, ZN => n2616);
   U2187 : OAI221_X1 port map( B1 => n2091, B2 => n2619, C1 => n2223, C2 => 
                           n2620, A => n2621, ZN => n2606);
   U2188 : AOI22_X1 port map( A1 => n2622, A2 => n3291, B1 => n2623, B2 => 
                           n3283, ZN => n2621);
   U2189 : OAI221_X1 port map( B1 => n2099, B2 => n2624, C1 => n2214, C2 => 
                           n2625, A => n2626, ZN => n2605);
   U2190 : AOI22_X1 port map( A1 => n2627, A2 => n3339, B1 => n2628, B2 => 
                           n3331, ZN => n2626);
   U2191 : AOI22_X1 port map( A1 => n2629, A2 => n3523, B1 => n2630, B2 => 
                           n2240, ZN => n2573);
   U2192 : OAI21_X1 port map( B1 => n2572, B2 => n2328, A => n2374, ZN => n1473
                           );
   U2193 : OAI211_X1 port map( C1 => n2572, C2 => n2353, A => n2631, B => n2632
                           , ZN => n1472);
   U2194 : AOI221_X1 port map( B1 => n2575, B2 => n3524, C1 => n2576, C2 => 
                           n2232, A => n2633, ZN => n2632);
   U2195 : AOI21_X1 port map( B1 => n2634, B2 => n2635, A => n2580, ZN => n2633
                           );
   U2196 : NOR4_X1 port map( A1 => n2636, A2 => n2637, A3 => n2638, A4 => n2639
                           , ZN => n2635);
   U2197 : OAI221_X1 port map( B1 => n2133, B2 => n2585, C1 => n2249, C2 => 
                           n2586, A => n2640, ZN => n2639);
   U2198 : AOI22_X1 port map( A1 => n2588, A2 => n3404, B1 => n2589, B2 => 
                           n3412, ZN => n2640);
   U2199 : OAI221_X1 port map( B1 => n2134, B2 => n2590, C1 => n2257, C2 => 
                           n2591, A => n2641, ZN => n2638);
   U2200 : AOI22_X1 port map( A1 => n2593, A2 => n3468, B1 => n2594, B2 => 
                           n3476, ZN => n2641);
   U2201 : OAI221_X1 port map( B1 => n2109, B2 => n2595, C1 => n2200, C2 => 
                           n2596, A => n2642, ZN => n2637);
   U2202 : AOI22_X1 port map( A1 => n2598, A2 => n2084, B1 => n2599, B2 => 
                           n2191, ZN => n2642);
   U2203 : OAI221_X1 port map( B1 => n2110, B2 => n2600, C1 => n2201, C2 => 
                           n2601, A => n2643, ZN => n2636);
   U2204 : AOI22_X1 port map( A1 => n2603, A2 => n3372, B1 => n2604, B2 => 
                           n3380, ZN => n2643);
   U2205 : NOR4_X1 port map( A1 => n2644, A2 => n2645, A3 => n2646, A4 => n2647
                           , ZN => n2634);
   U2206 : OAI221_X1 port map( B1 => n2124, B2 => n2609, C1 => n2273, C2 => 
                           n2610, A => n2648, ZN => n2647);
   U2207 : AOI22_X1 port map( A1 => n2612, A2 => n3428, B1 => n2613, B2 => 
                           n3420, ZN => n2648);
   U2208 : OAI221_X1 port map( B1 => n2148, B2 => n2614, C1 => n2265, C2 => 
                           n2615, A => n2649, ZN => n2646);
   U2209 : AOI22_X1 port map( A1 => n2617, A2 => n3492, B1 => n2618, B2 => 
                           n3484, ZN => n2649);
   U2210 : OAI221_X1 port map( B1 => n2092, B2 => n2619, C1 => n2224, C2 => 
                           n2620, A => n2650, ZN => n2645);
   U2211 : AOI22_X1 port map( A1 => n2622, A2 => n3284, B1 => n2623, B2 => 
                           n3276, ZN => n2650);
   U2212 : OAI221_X1 port map( B1 => n2100, B2 => n2624, C1 => n2215, C2 => 
                           n2625, A => n2651, ZN => n2644);
   U2213 : AOI22_X1 port map( A1 => n2627, A2 => n3332, B1 => n2628, B2 => 
                           n3324, ZN => n2651);
   U2214 : AOI22_X1 port map( A1 => n2629, A2 => n3516, B1 => n2630, B2 => 
                           n2241, ZN => n2631);
   U2215 : OAI21_X1 port map( B1 => n2572, B2 => n2329, A => n2374, ZN => n1471
                           );
   U2216 : OAI211_X1 port map( C1 => n2572, C2 => n2354, A => n2652, B => n2653
                           , ZN => n1470);
   U2217 : AOI221_X1 port map( B1 => n2575, B2 => n3530, C1 => n2576, C2 => 
                           n2233, A => n2654, ZN => n2653);
   U2218 : AOI21_X1 port map( B1 => n2655, B2 => n2656, A => n2580, ZN => n2654
                           );
   U2219 : NOR4_X1 port map( A1 => n2657, A2 => n2658, A3 => n2659, A4 => n2660
                           , ZN => n2656);
   U2220 : OAI221_X1 port map( B1 => n2135, B2 => n2585, C1 => n2250, C2 => 
                           n2586, A => n2661, ZN => n2660);
   U2221 : AOI22_X1 port map( A1 => n2588, A2 => n3410, B1 => n2589, B2 => 
                           n3418, ZN => n2661);
   U2222 : OAI221_X1 port map( B1 => n2136, B2 => n2590, C1 => n2258, C2 => 
                           n2591, A => n2662, ZN => n2659);
   U2223 : AOI22_X1 port map( A1 => n2593, A2 => n3474, B1 => n2594, B2 => 
                           n3482, ZN => n2662);
   U2224 : OAI221_X1 port map( B1 => n2111, B2 => n2595, C1 => n2202, C2 => 
                           n2596, A => n2663, ZN => n2658);
   U2225 : AOI22_X1 port map( A1 => n2598, A2 => n2085, B1 => n2599, B2 => 
                           n2192, ZN => n2663);
   U2226 : OAI221_X1 port map( B1 => n2112, B2 => n2600, C1 => n2203, C2 => 
                           n2601, A => n2664, ZN => n2657);
   U2227 : AOI22_X1 port map( A1 => n2603, A2 => n3378, B1 => n2604, B2 => 
                           n3386, ZN => n2664);
   U2228 : NOR4_X1 port map( A1 => n2665, A2 => n2666, A3 => n2667, A4 => n2668
                           , ZN => n2655);
   U2229 : OAI221_X1 port map( B1 => n2125, B2 => n2609, C1 => n2274, C2 => 
                           n2610, A => n2669, ZN => n2668);
   U2230 : AOI22_X1 port map( A1 => n2612, A2 => n3434, B1 => n2613, B2 => 
                           n3426, ZN => n2669);
   U2231 : OAI221_X1 port map( B1 => n2149, B2 => n2614, C1 => n2266, C2 => 
                           n2615, A => n2670, ZN => n2667);
   U2232 : AOI22_X1 port map( A1 => n2617, A2 => n3498, B1 => n2618, B2 => 
                           n3490, ZN => n2670);
   U2233 : OAI221_X1 port map( B1 => n2093, B2 => n2619, C1 => n2225, C2 => 
                           n2620, A => n2671, ZN => n2666);
   U2234 : AOI22_X1 port map( A1 => n2622, A2 => n3290, B1 => n2623, B2 => 
                           n3282, ZN => n2671);
   U2235 : OAI221_X1 port map( B1 => n2101, B2 => n2624, C1 => n2216, C2 => 
                           n2625, A => n2672, ZN => n2665);
   U2236 : AOI22_X1 port map( A1 => n2627, A2 => n3338, B1 => n2628, B2 => 
                           n3330, ZN => n2672);
   U2237 : AOI22_X1 port map( A1 => n2629, A2 => n3522, B1 => n2630, B2 => 
                           n2242, ZN => n2652);
   U2238 : OAI21_X1 port map( B1 => n2572, B2 => n2330, A => n2374, ZN => n1469
                           );
   U2239 : OAI211_X1 port map( C1 => n2572, C2 => n2355, A => n2673, B => n2674
                           , ZN => n1468);
   U2240 : AOI221_X1 port map( B1 => n2575, B2 => n3525, C1 => n2576, C2 => 
                           n2234, A => n2675, ZN => n2674);
   U2241 : AOI21_X1 port map( B1 => n2676, B2 => n2677, A => n2580, ZN => n2675
                           );
   U2242 : NOR4_X1 port map( A1 => n2678, A2 => n2679, A3 => n2680, A4 => n2681
                           , ZN => n2677);
   U2243 : OAI221_X1 port map( B1 => n2137, B2 => n2585, C1 => n2251, C2 => 
                           n2586, A => n2682, ZN => n2681);
   U2244 : AOI22_X1 port map( A1 => n2588, A2 => n3405, B1 => n2589, B2 => 
                           n3413, ZN => n2682);
   U2245 : OAI221_X1 port map( B1 => n2138, B2 => n2590, C1 => n2259, C2 => 
                           n2591, A => n2683, ZN => n2680);
   U2246 : AOI22_X1 port map( A1 => n2593, A2 => n3469, B1 => n2594, B2 => 
                           n3477, ZN => n2683);
   U2247 : OAI221_X1 port map( B1 => n2113, B2 => n2595, C1 => n2204, C2 => 
                           n2596, A => n2684, ZN => n2679);
   U2248 : AOI22_X1 port map( A1 => n2598, A2 => n2086, B1 => n2599, B2 => 
                           n2193, ZN => n2684);
   U2249 : OAI221_X1 port map( B1 => n2114, B2 => n2600, C1 => n2205, C2 => 
                           n2601, A => n2685, ZN => n2678);
   U2250 : AOI22_X1 port map( A1 => n2603, A2 => n3373, B1 => n2604, B2 => 
                           n3381, ZN => n2685);
   U2251 : NOR4_X1 port map( A1 => n2686, A2 => n2687, A3 => n2688, A4 => n2689
                           , ZN => n2676);
   U2252 : OAI221_X1 port map( B1 => n2126, B2 => n2609, C1 => n2275, C2 => 
                           n2610, A => n2690, ZN => n2689);
   U2253 : AOI22_X1 port map( A1 => n2612, A2 => n3429, B1 => n2613, B2 => 
                           n3421, ZN => n2690);
   U2254 : OAI221_X1 port map( B1 => n2150, B2 => n2614, C1 => n2267, C2 => 
                           n2615, A => n2691, ZN => n2688);
   U2255 : AOI22_X1 port map( A1 => n2617, A2 => n3493, B1 => n2618, B2 => 
                           n3485, ZN => n2691);
   U2256 : OAI221_X1 port map( B1 => n2094, B2 => n2619, C1 => n2226, C2 => 
                           n2620, A => n2692, ZN => n2687);
   U2257 : AOI22_X1 port map( A1 => n2622, A2 => n3285, B1 => n2623, B2 => 
                           n3277, ZN => n2692);
   U2258 : OAI221_X1 port map( B1 => n2102, B2 => n2624, C1 => n2217, C2 => 
                           n2625, A => n2693, ZN => n2686);
   U2259 : AOI22_X1 port map( A1 => n2627, A2 => n3333, B1 => n2628, B2 => 
                           n3325, ZN => n2693);
   U2260 : AOI22_X1 port map( A1 => n2629, A2 => n3517, B1 => n2630, B2 => 
                           n2243, ZN => n2673);
   U2261 : OAI21_X1 port map( B1 => n2572, B2 => n2331, A => n2374, ZN => n1467
                           );
   U2262 : OAI211_X1 port map( C1 => n2572, C2 => n2356, A => n2694, B => n2695
                           , ZN => n1466);
   U2263 : AOI221_X1 port map( B1 => n2575, B2 => n3529, C1 => n2576, C2 => 
                           n2235, A => n2696, ZN => n2695);
   U2264 : AOI21_X1 port map( B1 => n2697, B2 => n2698, A => n2580, ZN => n2696
                           );
   U2265 : NOR4_X1 port map( A1 => n2699, A2 => n2700, A3 => n2701, A4 => n2702
                           , ZN => n2698);
   U2266 : OAI221_X1 port map( B1 => n2139, B2 => n2585, C1 => n2252, C2 => 
                           n2586, A => n2703, ZN => n2702);
   U2267 : AOI22_X1 port map( A1 => n2588, A2 => n3409, B1 => n2589, B2 => 
                           n3417, ZN => n2703);
   U2268 : OAI221_X1 port map( B1 => n2140, B2 => n2590, C1 => n2260, C2 => 
                           n2591, A => n2704, ZN => n2701);
   U2269 : AOI22_X1 port map( A1 => n2593, A2 => n3473, B1 => n2594, B2 => 
                           n3481, ZN => n2704);
   U2270 : OAI221_X1 port map( B1 => n2115, B2 => n2595, C1 => n2206, C2 => 
                           n2596, A => n2705, ZN => n2700);
   U2271 : AOI22_X1 port map( A1 => n2598, A2 => n2087, B1 => n2599, B2 => 
                           n2194, ZN => n2705);
   U2272 : OAI221_X1 port map( B1 => n2116, B2 => n2600, C1 => n2207, C2 => 
                           n2601, A => n2706, ZN => n2699);
   U2273 : AOI22_X1 port map( A1 => n2603, A2 => n3377, B1 => n2604, B2 => 
                           n3385, ZN => n2706);
   U2274 : NOR4_X1 port map( A1 => n2707, A2 => n2708, A3 => n2709, A4 => n2710
                           , ZN => n2697);
   U2275 : OAI221_X1 port map( B1 => n2127, B2 => n2609, C1 => n2276, C2 => 
                           n2610, A => n2711, ZN => n2710);
   U2276 : AOI22_X1 port map( A1 => n2612, A2 => n3433, B1 => n2613, B2 => 
                           n3425, ZN => n2711);
   U2277 : OAI221_X1 port map( B1 => n2151, B2 => n2614, C1 => n2268, C2 => 
                           n2615, A => n2712, ZN => n2709);
   U2278 : AOI22_X1 port map( A1 => n2617, A2 => n3497, B1 => n2618, B2 => 
                           n3489, ZN => n2712);
   U2279 : OAI221_X1 port map( B1 => n2095, B2 => n2619, C1 => n2227, C2 => 
                           n2620, A => n2713, ZN => n2708);
   U2280 : AOI22_X1 port map( A1 => n2622, A2 => n3289, B1 => n2623, B2 => 
                           n3281, ZN => n2713);
   U2281 : OAI221_X1 port map( B1 => n2103, B2 => n2624, C1 => n2218, C2 => 
                           n2625, A => n2714, ZN => n2707);
   U2282 : AOI22_X1 port map( A1 => n2627, A2 => n3337, B1 => n2628, B2 => 
                           n3329, ZN => n2714);
   U2283 : AOI22_X1 port map( A1 => n2629, A2 => n3521, B1 => n2630, B2 => 
                           n2244, ZN => n2694);
   U2284 : OAI21_X1 port map( B1 => n2572, B2 => n2332, A => n2374, ZN => n1465
                           );
   U2285 : OAI211_X1 port map( C1 => n2572, C2 => n2357, A => n2715, B => n2716
                           , ZN => n1464);
   U2286 : AOI221_X1 port map( B1 => n2575, B2 => n3526, C1 => n2576, C2 => 
                           n2236, A => n2717, ZN => n2716);
   U2287 : AOI21_X1 port map( B1 => n2718, B2 => n2719, A => n2580, ZN => n2717
                           );
   U2288 : NOR4_X1 port map( A1 => n2720, A2 => n2721, A3 => n2722, A4 => n2723
                           , ZN => n2719);
   U2289 : OAI221_X1 port map( B1 => n2141, B2 => n2585, C1 => n2253, C2 => 
                           n2586, A => n2724, ZN => n2723);
   U2290 : AOI22_X1 port map( A1 => n2588, A2 => n3406, B1 => n2589, B2 => 
                           n3414, ZN => n2724);
   U2291 : OAI221_X1 port map( B1 => n2142, B2 => n2590, C1 => n2261, C2 => 
                           n2591, A => n2725, ZN => n2722);
   U2292 : AOI22_X1 port map( A1 => n2593, A2 => n3470, B1 => n2594, B2 => 
                           n3478, ZN => n2725);
   U2293 : OAI221_X1 port map( B1 => n2117, B2 => n2595, C1 => n2208, C2 => 
                           n2596, A => n2726, ZN => n2721);
   U2294 : AOI22_X1 port map( A1 => n2598, A2 => n2088, B1 => n2599, B2 => 
                           n2195, ZN => n2726);
   U2295 : OAI221_X1 port map( B1 => n2118, B2 => n2600, C1 => n2209, C2 => 
                           n2601, A => n2727, ZN => n2720);
   U2296 : AOI22_X1 port map( A1 => n2603, A2 => n3374, B1 => n2604, B2 => 
                           n3382, ZN => n2727);
   U2297 : NOR4_X1 port map( A1 => n2728, A2 => n2729, A3 => n2730, A4 => n2731
                           , ZN => n2718);
   U2298 : OAI221_X1 port map( B1 => n2128, B2 => n2609, C1 => n2277, C2 => 
                           n2610, A => n2732, ZN => n2731);
   U2299 : AOI22_X1 port map( A1 => n2612, A2 => n3430, B1 => n2613, B2 => 
                           n3422, ZN => n2732);
   U2300 : OAI221_X1 port map( B1 => n2152, B2 => n2614, C1 => n2269, C2 => 
                           n2615, A => n2733, ZN => n2730);
   U2301 : AOI22_X1 port map( A1 => n2617, A2 => n3494, B1 => n2618, B2 => 
                           n3486, ZN => n2733);
   U2302 : OAI221_X1 port map( B1 => n2096, B2 => n2619, C1 => n2228, C2 => 
                           n2620, A => n2734, ZN => n2729);
   U2303 : AOI22_X1 port map( A1 => n2622, A2 => n3286, B1 => n2623, B2 => 
                           n3278, ZN => n2734);
   U2304 : OAI221_X1 port map( B1 => n2104, B2 => n2624, C1 => n2219, C2 => 
                           n2625, A => n2735, ZN => n2728);
   U2305 : AOI22_X1 port map( A1 => n2627, A2 => n3334, B1 => n2628, B2 => 
                           n3326, ZN => n2735);
   U2306 : AOI22_X1 port map( A1 => n2629, A2 => n3518, B1 => n2630, B2 => 
                           n2245, ZN => n2715);
   U2307 : OAI21_X1 port map( B1 => n2572, B2 => n2333, A => n2374, ZN => n1463
                           );
   U2308 : OAI211_X1 port map( C1 => n2572, C2 => n2358, A => n2736, B => n2737
                           , ZN => n1462);
   U2309 : AOI221_X1 port map( B1 => n2575, B2 => n3528, C1 => n2576, C2 => 
                           n2237, A => n2738, ZN => n2737);
   U2310 : AOI21_X1 port map( B1 => n2739, B2 => n2740, A => n2580, ZN => n2738
                           );
   U2311 : NOR4_X1 port map( A1 => n2741, A2 => n2742, A3 => n2743, A4 => n2744
                           , ZN => n2740);
   U2312 : OAI221_X1 port map( B1 => n2143, B2 => n2585, C1 => n2254, C2 => 
                           n2586, A => n2745, ZN => n2744);
   U2313 : AOI22_X1 port map( A1 => n2588, A2 => n3408, B1 => n2589, B2 => 
                           n3416, ZN => n2745);
   U2314 : OAI221_X1 port map( B1 => n2144, B2 => n2590, C1 => n2262, C2 => 
                           n2591, A => n2746, ZN => n2743);
   U2315 : AOI22_X1 port map( A1 => n2593, A2 => n3472, B1 => n2594, B2 => 
                           n3480, ZN => n2746);
   U2316 : OAI221_X1 port map( B1 => n2119, B2 => n2595, C1 => n2210, C2 => 
                           n2596, A => n2747, ZN => n2742);
   U2317 : AOI22_X1 port map( A1 => n2598, A2 => n2089, B1 => n2599, B2 => 
                           n2196, ZN => n2747);
   U2318 : OAI221_X1 port map( B1 => n2120, B2 => n2600, C1 => n2211, C2 => 
                           n2601, A => n2748, ZN => n2741);
   U2319 : AOI22_X1 port map( A1 => n2603, A2 => n3376, B1 => n2604, B2 => 
                           n3384, ZN => n2748);
   U2320 : NOR4_X1 port map( A1 => n2749, A2 => n2750, A3 => n2751, A4 => n2752
                           , ZN => n2739);
   U2321 : OAI221_X1 port map( B1 => n2129, B2 => n2609, C1 => n2278, C2 => 
                           n2610, A => n2753, ZN => n2752);
   U2322 : AOI22_X1 port map( A1 => n2612, A2 => n3432, B1 => n2613, B2 => 
                           n3424, ZN => n2753);
   U2323 : OAI221_X1 port map( B1 => n2153, B2 => n2614, C1 => n2270, C2 => 
                           n2615, A => n2754, ZN => n2751);
   U2324 : AOI22_X1 port map( A1 => n2617, A2 => n3496, B1 => n2618, B2 => 
                           n3488, ZN => n2754);
   U2325 : OAI221_X1 port map( B1 => n2097, B2 => n2619, C1 => n2229, C2 => 
                           n2620, A => n2755, ZN => n2750);
   U2326 : AOI22_X1 port map( A1 => n2622, A2 => n3288, B1 => n2623, B2 => 
                           n3280, ZN => n2755);
   U2327 : OAI221_X1 port map( B1 => n2105, B2 => n2624, C1 => n2220, C2 => 
                           n2625, A => n2756, ZN => n2749);
   U2328 : AOI22_X1 port map( A1 => n2627, A2 => n3336, B1 => n2628, B2 => 
                           n3328, ZN => n2756);
   U2329 : AOI22_X1 port map( A1 => n2629, A2 => n3520, B1 => n2630, B2 => 
                           n2246, ZN => n2736);
   U2330 : OAI21_X1 port map( B1 => n2572, B2 => n2334, A => n2374, ZN => n1461
                           );
   U2331 : OAI211_X1 port map( C1 => n2572, C2 => n2359, A => n2757, B => n2758
                           , ZN => n1460);
   U2332 : AOI221_X1 port map( B1 => n2575, B2 => n3527, C1 => n2576, C2 => 
                           n2238, A => n2759, ZN => n2758);
   U2333 : AOI21_X1 port map( B1 => n2760, B2 => n2761, A => n2580, ZN => n2759
                           );
   U2334 : NAND2_X1 port map( A1 => n2762, A2 => n2572, ZN => n2580);
   U2335 : NOR4_X1 port map( A1 => n2763, A2 => n2764, A3 => n2765, A4 => n2766
                           , ZN => n2761);
   U2336 : OAI221_X1 port map( B1 => n2145, B2 => n2585, C1 => n2255, C2 => 
                           n2586, A => n2767, ZN => n2766);
   U2337 : AOI22_X1 port map( A1 => n2588, A2 => n3407, B1 => n2589, B2 => 
                           n3415, ZN => n2767);
   U2338 : AND2_X1 port map( A1 => n2768, A2 => n2769, ZN => n2589);
   U2339 : AND2_X1 port map( A1 => n2770, A2 => n2769, ZN => n2588);
   U2340 : NAND2_X1 port map( A1 => n2768, A2 => n2771, ZN => n2586);
   U2341 : NAND2_X1 port map( A1 => n2770, A2 => n2771, ZN => n2585);
   U2342 : OAI221_X1 port map( B1 => n2146, B2 => n2590, C1 => n2263, C2 => 
                           n2591, A => n2772, ZN => n2765);
   U2343 : AOI22_X1 port map( A1 => n2593, A2 => n3471, B1 => n2594, B2 => 
                           n3479, ZN => n2772);
   U2344 : AND2_X1 port map( A1 => n2773, A2 => n2769, ZN => n2594);
   U2345 : AND2_X1 port map( A1 => n2774, A2 => n2769, ZN => n2593);
   U2346 : NAND2_X1 port map( A1 => n2773, A2 => n2771, ZN => n2591);
   U2347 : NAND2_X1 port map( A1 => n2774, A2 => n2771, ZN => n2590);
   U2348 : OAI221_X1 port map( B1 => n2121, B2 => n2595, C1 => n2212, C2 => 
                           n2596, A => n2775, ZN => n2764);
   U2349 : AOI22_X1 port map( A1 => n2598, A2 => n2090, B1 => n2599, B2 => 
                           n2197, ZN => n2775);
   U2350 : AND2_X1 port map( A1 => n2776, A2 => n2777, ZN => n2599);
   U2351 : AND2_X1 port map( A1 => n2776, A2 => n2778, ZN => n2598);
   U2352 : NAND2_X1 port map( A1 => n2777, A2 => n2771, ZN => n2596);
   U2353 : NAND2_X1 port map( A1 => n2778, A2 => n2771, ZN => n2595);
   U2354 : OAI221_X1 port map( B1 => n2122, B2 => n2600, C1 => n2213, C2 => 
                           n2601, A => n2779, ZN => n2763);
   U2355 : AOI22_X1 port map( A1 => n2603, A2 => n3375, B1 => n2604, B2 => 
                           n3383, ZN => n2779);
   U2356 : AND2_X1 port map( A1 => n2771, A2 => n2780, ZN => n2604);
   U2357 : AND2_X1 port map( A1 => n2771, A2 => n2781, ZN => n2603);
   U2358 : NOR2_X1 port map( A1 => N108, A2 => N109, ZN => n2771);
   U2359 : NAND2_X1 port map( A1 => n2780, A2 => n2769, ZN => n2601);
   U2360 : NAND2_X1 port map( A1 => n2769, A2 => n2781, ZN => n2600);
   U2361 : NOR4_X1 port map( A1 => n2782, A2 => n2783, A3 => n2784, A4 => n2785
                           , ZN => n2760);
   U2362 : OAI221_X1 port map( B1 => n2130, B2 => n2609, C1 => n2279, C2 => 
                           n2610, A => n2786, ZN => n2785);
   U2363 : AOI22_X1 port map( A1 => n2612, A2 => n3431, B1 => n2613, B2 => 
                           n3423, ZN => n2786);
   U2364 : AND2_X1 port map( A1 => n2787, A2 => n2770, ZN => n2613);
   U2365 : AND2_X1 port map( A1 => n2787, A2 => n2768, ZN => n2612);
   U2366 : NAND2_X1 port map( A1 => n2770, A2 => n2776, ZN => n2610);
   U2367 : NOR3_X1 port map( A1 => n2788, A2 => N111, A3 => n2789, ZN => n2770)
                           ;
   U2368 : NAND2_X1 port map( A1 => n2768, A2 => n2776, ZN => n2609);
   U2369 : NOR3_X1 port map( A1 => N107, A2 => N111, A3 => n2789, ZN => n2768);
   U2370 : OAI221_X1 port map( B1 => n2154, B2 => n2614, C1 => n2271, C2 => 
                           n2615, A => n2790, ZN => n2784);
   U2371 : AOI22_X1 port map( A1 => n2617, A2 => n3495, B1 => n2618, B2 => 
                           n3487, ZN => n2790);
   U2372 : AND2_X1 port map( A1 => n2787, A2 => n2774, ZN => n2618);
   U2373 : AND2_X1 port map( A1 => n2787, A2 => n2773, ZN => n2617);
   U2374 : NAND2_X1 port map( A1 => n2774, A2 => n2776, ZN => n2615);
   U2375 : NOR3_X1 port map( A1 => N110, A2 => N111, A3 => n2788, ZN => n2774);
   U2376 : NAND2_X1 port map( A1 => n2773, A2 => n2776, ZN => n2614);
   U2377 : NOR3_X1 port map( A1 => N110, A2 => N111, A3 => N107, ZN => n2773);
   U2378 : OAI221_X1 port map( B1 => n2098, B2 => n2619, C1 => n2230, C2 => 
                           n2620, A => n2791, ZN => n2783);
   U2379 : AOI22_X1 port map( A1 => n2622, A2 => n3287, B1 => n2623, B2 => 
                           n3279, ZN => n2791);
   U2380 : AND2_X1 port map( A1 => n2778, A2 => n2769, ZN => n2623);
   U2381 : AND2_X1 port map( A1 => n2777, A2 => n2769, ZN => n2622);
   U2382 : NOR2_X1 port map( A1 => n2792, A2 => N108, ZN => n2769);
   U2383 : NAND2_X1 port map( A1 => n2787, A2 => n2778, ZN => n2620);
   U2384 : NOR3_X1 port map( A1 => n2793, A2 => n2788, A3 => n2789, ZN => n2778
                           );
   U2385 : NAND2_X1 port map( A1 => n2787, A2 => n2777, ZN => n2619);
   U2386 : NOR3_X1 port map( A1 => n2793, A2 => N107, A3 => n2789, ZN => n2777)
                           ;
   U2387 : INV_X1 port map( A => N110, ZN => n2789);
   U2388 : OAI221_X1 port map( B1 => n2106, B2 => n2624, C1 => n2221, C2 => 
                           n2625, A => n2794, ZN => n2782);
   U2389 : AOI22_X1 port map( A1 => n2627, A2 => n3335, B1 => n2628, B2 => 
                           n3327, ZN => n2794);
   U2390 : AND2_X1 port map( A1 => n2776, A2 => n2781, ZN => n2628);
   U2391 : AND2_X1 port map( A1 => n2776, A2 => n2780, ZN => n2627);
   U2392 : NOR2_X1 port map( A1 => n2795, A2 => n2792, ZN => n2776);
   U2393 : INV_X1 port map( A => N109, ZN => n2792);
   U2394 : NAND2_X1 port map( A1 => n2787, A2 => n2781, ZN => n2625);
   U2395 : NOR3_X1 port map( A1 => n2788, A2 => N110, A3 => n2793, ZN => n2781)
                           ;
   U2396 : INV_X1 port map( A => N107, ZN => n2788);
   U2397 : NAND2_X1 port map( A1 => n2787, A2 => n2780, ZN => n2624);
   U2398 : NOR3_X1 port map( A1 => N107, A2 => N110, A3 => n2793, ZN => n2780);
   U2399 : INV_X1 port map( A => N111, ZN => n2793);
   U2400 : NOR2_X1 port map( A1 => n2795, A2 => N109, ZN => n2787);
   U2401 : INV_X1 port map( A => N108, ZN => n2795);
   U2402 : AND3_X1 port map( A1 => n2796, A2 => n2797, A3 => n2798, ZN => n2576
                           );
   U2403 : AND3_X1 port map( A1 => n2798, A2 => n2796, A3 => ADD_RD1(1), ZN => 
                           n2575);
   U2404 : INV_X1 port map( A => ADD_RD1(0), ZN => n2796);
   U2405 : AOI22_X1 port map( A1 => n2629, A2 => n3519, B1 => n2630, B2 => 
                           n2247, ZN => n2757);
   U2406 : AND3_X1 port map( A1 => n2798, A2 => n2797, A3 => ADD_RD1(0), ZN => 
                           n2630);
   U2407 : INV_X1 port map( A => ADD_RD1(1), ZN => n2797);
   U2408 : AND3_X1 port map( A1 => ADD_RD1(1), A2 => n2798, A3 => ADD_RD1(0), 
                           ZN => n2629);
   U2409 : AND2_X1 port map( A1 => n2799, A2 => n2572, ZN => n2798);
   U2410 : OAI21_X1 port map( B1 => n2572, B2 => n2335, A => n2374, ZN => n1459
                           );
   U2411 : NAND2_X1 port map( A1 => n2800, A2 => n2374, ZN => n2572);
   U2412 : NAND2_X1 port map( A1 => RD1, A2 => n2432, ZN => n2800);
   U2413 : OAI211_X1 port map( C1 => n2801, C2 => n2360, A => n2802, B => n2803
                           , ZN => n1458);
   U2414 : AOI221_X1 port map( B1 => n2804, B2 => n3531, C1 => n2805, C2 => 
                           n2231, A => n2806, ZN => n2803);
   U2415 : AOI21_X1 port map( B1 => n2807, B2 => n2808, A => n2809, ZN => n2806
                           );
   U2416 : NOR4_X1 port map( A1 => n2810, A2 => n2811, A3 => n2812, A4 => n2813
                           , ZN => n2808);
   U2417 : OAI221_X1 port map( B1 => n2131, B2 => n2814, C1 => n2248, C2 => 
                           n2815, A => n2816, ZN => n2813);
   U2418 : AOI22_X1 port map( A1 => n2817, A2 => n3411, B1 => n2818, B2 => 
                           n3419, ZN => n2816);
   U2419 : OAI221_X1 port map( B1 => n2132, B2 => n2819, C1 => n2256, C2 => 
                           n2820, A => n2821, ZN => n2812);
   U2420 : AOI22_X1 port map( A1 => n2822, A2 => n3475, B1 => n2823, B2 => 
                           n3483, ZN => n2821);
   U2421 : OAI221_X1 port map( B1 => n2107, B2 => n2824, C1 => n2198, C2 => 
                           n2825, A => n2826, ZN => n2811);
   U2422 : AOI22_X1 port map( A1 => n2827, A2 => n2083, B1 => n2828, B2 => 
                           n2190, ZN => n2826);
   U2423 : OAI221_X1 port map( B1 => n2108, B2 => n2829, C1 => n2199, C2 => 
                           n2830, A => n2831, ZN => n2810);
   U2424 : AOI22_X1 port map( A1 => n2832, A2 => n3379, B1 => n2833, B2 => 
                           n3387, ZN => n2831);
   U2425 : NOR4_X1 port map( A1 => n2834, A2 => n2835, A3 => n2836, A4 => n2837
                           , ZN => n2807);
   U2426 : OAI221_X1 port map( B1 => n2123, B2 => n2838, C1 => n2272, C2 => 
                           n2839, A => n2840, ZN => n2837);
   U2427 : AOI22_X1 port map( A1 => n2841, A2 => n3435, B1 => n2842, B2 => 
                           n3427, ZN => n2840);
   U2428 : OAI221_X1 port map( B1 => n2147, B2 => n2843, C1 => n2264, C2 => 
                           n2844, A => n2845, ZN => n2836);
   U2429 : AOI22_X1 port map( A1 => n2846, A2 => n3499, B1 => n2847, B2 => 
                           n3491, ZN => n2845);
   U2430 : OAI221_X1 port map( B1 => n2091, B2 => n2848, C1 => n2223, C2 => 
                           n2849, A => n2850, ZN => n2835);
   U2431 : AOI22_X1 port map( A1 => n2851, A2 => n3291, B1 => n2852, B2 => 
                           n3283, ZN => n2850);
   U2432 : OAI221_X1 port map( B1 => n2099, B2 => n2853, C1 => n2214, C2 => 
                           n2854, A => n2855, ZN => n2834);
   U2433 : AOI22_X1 port map( A1 => n2856, A2 => n3339, B1 => n2857, B2 => 
                           n3331, ZN => n2855);
   U2434 : AOI22_X1 port map( A1 => n2858, A2 => n3523, B1 => n2859, B2 => 
                           n2240, ZN => n2802);
   U2435 : OAI21_X1 port map( B1 => n2801, B2 => n2336, A => n2374, ZN => n1457
                           );
   U2436 : OAI211_X1 port map( C1 => n2801, C2 => n2361, A => n2860, B => n2861
                           , ZN => n1456);
   U2437 : AOI221_X1 port map( B1 => n2804, B2 => n3524, C1 => n2805, C2 => 
                           n2232, A => n2862, ZN => n2861);
   U2438 : AOI21_X1 port map( B1 => n2863, B2 => n2864, A => n2809, ZN => n2862
                           );
   U2439 : NOR4_X1 port map( A1 => n2865, A2 => n2866, A3 => n2867, A4 => n2868
                           , ZN => n2864);
   U2440 : OAI221_X1 port map( B1 => n2133, B2 => n2814, C1 => n2249, C2 => 
                           n2815, A => n2869, ZN => n2868);
   U2441 : AOI22_X1 port map( A1 => n2817, A2 => n3404, B1 => n2818, B2 => 
                           n3412, ZN => n2869);
   U2442 : OAI221_X1 port map( B1 => n2134, B2 => n2819, C1 => n2257, C2 => 
                           n2820, A => n2870, ZN => n2867);
   U2443 : AOI22_X1 port map( A1 => n2822, A2 => n3468, B1 => n2823, B2 => 
                           n3476, ZN => n2870);
   U2444 : OAI221_X1 port map( B1 => n2109, B2 => n2824, C1 => n2200, C2 => 
                           n2825, A => n2871, ZN => n2866);
   U2445 : AOI22_X1 port map( A1 => n2827, A2 => n2084, B1 => n2828, B2 => 
                           n2191, ZN => n2871);
   U2446 : OAI221_X1 port map( B1 => n2110, B2 => n2829, C1 => n2201, C2 => 
                           n2830, A => n2872, ZN => n2865);
   U2447 : AOI22_X1 port map( A1 => n2832, A2 => n3372, B1 => n2833, B2 => 
                           n3380, ZN => n2872);
   U2448 : NOR4_X1 port map( A1 => n2873, A2 => n2874, A3 => n2875, A4 => n2876
                           , ZN => n2863);
   U2449 : OAI221_X1 port map( B1 => n2124, B2 => n2838, C1 => n2273, C2 => 
                           n2839, A => n2877, ZN => n2876);
   U2450 : AOI22_X1 port map( A1 => n2841, A2 => n3428, B1 => n2842, B2 => 
                           n3420, ZN => n2877);
   U2451 : OAI221_X1 port map( B1 => n2148, B2 => n2843, C1 => n2265, C2 => 
                           n2844, A => n2878, ZN => n2875);
   U2452 : AOI22_X1 port map( A1 => n2846, A2 => n3492, B1 => n2847, B2 => 
                           n3484, ZN => n2878);
   U2453 : OAI221_X1 port map( B1 => n2092, B2 => n2848, C1 => n2224, C2 => 
                           n2849, A => n2879, ZN => n2874);
   U2454 : AOI22_X1 port map( A1 => n2851, A2 => n3284, B1 => n2852, B2 => 
                           n3276, ZN => n2879);
   U2455 : OAI221_X1 port map( B1 => n2100, B2 => n2853, C1 => n2215, C2 => 
                           n2854, A => n2880, ZN => n2873);
   U2456 : AOI22_X1 port map( A1 => n2856, A2 => n3332, B1 => n2857, B2 => 
                           n3324, ZN => n2880);
   U2457 : AOI22_X1 port map( A1 => n2858, A2 => n3516, B1 => n2859, B2 => 
                           n2241, ZN => n2860);
   U2458 : OAI21_X1 port map( B1 => n2801, B2 => n2337, A => n2374, ZN => n1455
                           );
   U2459 : OAI211_X1 port map( C1 => n2801, C2 => n2362, A => n2881, B => n2882
                           , ZN => n1454);
   U2460 : AOI221_X1 port map( B1 => n2804, B2 => n3530, C1 => n2805, C2 => 
                           n2233, A => n2883, ZN => n2882);
   U2461 : AOI21_X1 port map( B1 => n2884, B2 => n2885, A => n2809, ZN => n2883
                           );
   U2462 : NOR4_X1 port map( A1 => n2886, A2 => n2887, A3 => n2888, A4 => n2889
                           , ZN => n2885);
   U2463 : OAI221_X1 port map( B1 => n2135, B2 => n2814, C1 => n2250, C2 => 
                           n2815, A => n2890, ZN => n2889);
   U2464 : AOI22_X1 port map( A1 => n2817, A2 => n3410, B1 => n2818, B2 => 
                           n3418, ZN => n2890);
   U2465 : OAI221_X1 port map( B1 => n2136, B2 => n2819, C1 => n2258, C2 => 
                           n2820, A => n2891, ZN => n2888);
   U2466 : AOI22_X1 port map( A1 => n2822, A2 => n3474, B1 => n2823, B2 => 
                           n3482, ZN => n2891);
   U2467 : OAI221_X1 port map( B1 => n2111, B2 => n2824, C1 => n2202, C2 => 
                           n2825, A => n2892, ZN => n2887);
   U2468 : AOI22_X1 port map( A1 => n2827, A2 => n2085, B1 => n2828, B2 => 
                           n2192, ZN => n2892);
   U2469 : OAI221_X1 port map( B1 => n2112, B2 => n2829, C1 => n2203, C2 => 
                           n2830, A => n2893, ZN => n2886);
   U2470 : AOI22_X1 port map( A1 => n2832, A2 => n3378, B1 => n2833, B2 => 
                           n3386, ZN => n2893);
   U2471 : NOR4_X1 port map( A1 => n2894, A2 => n2895, A3 => n2896, A4 => n2897
                           , ZN => n2884);
   U2472 : OAI221_X1 port map( B1 => n2125, B2 => n2838, C1 => n2274, C2 => 
                           n2839, A => n2898, ZN => n2897);
   U2473 : AOI22_X1 port map( A1 => n2841, A2 => n3434, B1 => n2842, B2 => 
                           n3426, ZN => n2898);
   U2474 : OAI221_X1 port map( B1 => n2149, B2 => n2843, C1 => n2266, C2 => 
                           n2844, A => n2899, ZN => n2896);
   U2475 : AOI22_X1 port map( A1 => n2846, A2 => n3498, B1 => n2847, B2 => 
                           n3490, ZN => n2899);
   U2476 : OAI221_X1 port map( B1 => n2093, B2 => n2848, C1 => n2225, C2 => 
                           n2849, A => n2900, ZN => n2895);
   U2477 : AOI22_X1 port map( A1 => n2851, A2 => n3290, B1 => n2852, B2 => 
                           n3282, ZN => n2900);
   U2478 : OAI221_X1 port map( B1 => n2101, B2 => n2853, C1 => n2216, C2 => 
                           n2854, A => n2901, ZN => n2894);
   U2479 : AOI22_X1 port map( A1 => n2856, A2 => n3338, B1 => n2857, B2 => 
                           n3330, ZN => n2901);
   U2480 : AOI22_X1 port map( A1 => n2858, A2 => n3522, B1 => n2859, B2 => 
                           n2242, ZN => n2881);
   U2481 : OAI21_X1 port map( B1 => n2801, B2 => n2338, A => n2374, ZN => n1453
                           );
   U2482 : OAI211_X1 port map( C1 => n2801, C2 => n2363, A => n2902, B => n2903
                           , ZN => n1452);
   U2483 : AOI221_X1 port map( B1 => n2804, B2 => n3525, C1 => n2805, C2 => 
                           n2234, A => n2904, ZN => n2903);
   U2484 : AOI21_X1 port map( B1 => n2905, B2 => n2906, A => n2809, ZN => n2904
                           );
   U2485 : NOR4_X1 port map( A1 => n2907, A2 => n2908, A3 => n2909, A4 => n2910
                           , ZN => n2906);
   U2486 : OAI221_X1 port map( B1 => n2137, B2 => n2814, C1 => n2251, C2 => 
                           n2815, A => n2911, ZN => n2910);
   U2487 : AOI22_X1 port map( A1 => n2817, A2 => n3405, B1 => n2818, B2 => 
                           n3413, ZN => n2911);
   U2488 : OAI221_X1 port map( B1 => n2138, B2 => n2819, C1 => n2259, C2 => 
                           n2820, A => n2912, ZN => n2909);
   U2489 : AOI22_X1 port map( A1 => n2822, A2 => n3469, B1 => n2823, B2 => 
                           n3477, ZN => n2912);
   U2490 : OAI221_X1 port map( B1 => n2113, B2 => n2824, C1 => n2204, C2 => 
                           n2825, A => n2913, ZN => n2908);
   U2491 : AOI22_X1 port map( A1 => n2827, A2 => n2086, B1 => n2828, B2 => 
                           n2193, ZN => n2913);
   U2492 : OAI221_X1 port map( B1 => n2114, B2 => n2829, C1 => n2205, C2 => 
                           n2830, A => n2914, ZN => n2907);
   U2493 : AOI22_X1 port map( A1 => n2832, A2 => n3373, B1 => n2833, B2 => 
                           n3381, ZN => n2914);
   U2494 : NOR4_X1 port map( A1 => n2915, A2 => n2916, A3 => n2917, A4 => n2918
                           , ZN => n2905);
   U2495 : OAI221_X1 port map( B1 => n2126, B2 => n2838, C1 => n2275, C2 => 
                           n2839, A => n2919, ZN => n2918);
   U2496 : AOI22_X1 port map( A1 => n2841, A2 => n3429, B1 => n2842, B2 => 
                           n3421, ZN => n2919);
   U2497 : OAI221_X1 port map( B1 => n2150, B2 => n2843, C1 => n2267, C2 => 
                           n2844, A => n2920, ZN => n2917);
   U2498 : AOI22_X1 port map( A1 => n2846, A2 => n3493, B1 => n2847, B2 => 
                           n3485, ZN => n2920);
   U2499 : OAI221_X1 port map( B1 => n2094, B2 => n2848, C1 => n2226, C2 => 
                           n2849, A => n2921, ZN => n2916);
   U2500 : AOI22_X1 port map( A1 => n2851, A2 => n3285, B1 => n2852, B2 => 
                           n3277, ZN => n2921);
   U2501 : OAI221_X1 port map( B1 => n2102, B2 => n2853, C1 => n2217, C2 => 
                           n2854, A => n2922, ZN => n2915);
   U2502 : AOI22_X1 port map( A1 => n2856, A2 => n3333, B1 => n2857, B2 => 
                           n3325, ZN => n2922);
   U2503 : AOI22_X1 port map( A1 => n2858, A2 => n3517, B1 => n2859, B2 => 
                           n2243, ZN => n2902);
   U2504 : OAI21_X1 port map( B1 => n2801, B2 => n2339, A => n2374, ZN => n1451
                           );
   U2505 : OAI211_X1 port map( C1 => n2801, C2 => n2364, A => n2923, B => n2924
                           , ZN => n1450);
   U2506 : AOI221_X1 port map( B1 => n2804, B2 => n3529, C1 => n2805, C2 => 
                           n2235, A => n2925, ZN => n2924);
   U2507 : AOI21_X1 port map( B1 => n2926, B2 => n2927, A => n2809, ZN => n2925
                           );
   U2508 : NOR4_X1 port map( A1 => n2928, A2 => n2929, A3 => n2930, A4 => n2931
                           , ZN => n2927);
   U2509 : OAI221_X1 port map( B1 => n2139, B2 => n2814, C1 => n2252, C2 => 
                           n2815, A => n2932, ZN => n2931);
   U2510 : AOI22_X1 port map( A1 => n2817, A2 => n3409, B1 => n2818, B2 => 
                           n3417, ZN => n2932);
   U2511 : OAI221_X1 port map( B1 => n2140, B2 => n2819, C1 => n2260, C2 => 
                           n2820, A => n2933, ZN => n2930);
   U2512 : AOI22_X1 port map( A1 => n2822, A2 => n3473, B1 => n2823, B2 => 
                           n3481, ZN => n2933);
   U2513 : OAI221_X1 port map( B1 => n2115, B2 => n2824, C1 => n2206, C2 => 
                           n2825, A => n2934, ZN => n2929);
   U2514 : AOI22_X1 port map( A1 => n2827, A2 => n2087, B1 => n2828, B2 => 
                           n2194, ZN => n2934);
   U2515 : OAI221_X1 port map( B1 => n2116, B2 => n2829, C1 => n2207, C2 => 
                           n2830, A => n2935, ZN => n2928);
   U2516 : AOI22_X1 port map( A1 => n2832, A2 => n3377, B1 => n2833, B2 => 
                           n3385, ZN => n2935);
   U2517 : NOR4_X1 port map( A1 => n2936, A2 => n2937, A3 => n2938, A4 => n2939
                           , ZN => n2926);
   U2518 : OAI221_X1 port map( B1 => n2127, B2 => n2838, C1 => n2276, C2 => 
                           n2839, A => n2940, ZN => n2939);
   U2519 : AOI22_X1 port map( A1 => n2841, A2 => n3433, B1 => n2842, B2 => 
                           n3425, ZN => n2940);
   U2520 : OAI221_X1 port map( B1 => n2151, B2 => n2843, C1 => n2268, C2 => 
                           n2844, A => n2941, ZN => n2938);
   U2521 : AOI22_X1 port map( A1 => n2846, A2 => n3497, B1 => n2847, B2 => 
                           n3489, ZN => n2941);
   U2522 : OAI221_X1 port map( B1 => n2095, B2 => n2848, C1 => n2227, C2 => 
                           n2849, A => n2942, ZN => n2937);
   U2523 : AOI22_X1 port map( A1 => n2851, A2 => n3289, B1 => n2852, B2 => 
                           n3281, ZN => n2942);
   U2524 : OAI221_X1 port map( B1 => n2103, B2 => n2853, C1 => n2218, C2 => 
                           n2854, A => n2943, ZN => n2936);
   U2525 : AOI22_X1 port map( A1 => n2856, A2 => n3337, B1 => n2857, B2 => 
                           n3329, ZN => n2943);
   U2526 : AOI22_X1 port map( A1 => n2858, A2 => n3521, B1 => n2859, B2 => 
                           n2244, ZN => n2923);
   U2527 : OAI21_X1 port map( B1 => n2801, B2 => n2340, A => n2374, ZN => n1449
                           );
   U2528 : OAI211_X1 port map( C1 => n2801, C2 => n2365, A => n2944, B => n2945
                           , ZN => n1448);
   U2529 : AOI221_X1 port map( B1 => n2804, B2 => n3526, C1 => n2805, C2 => 
                           n2236, A => n2946, ZN => n2945);
   U2530 : AOI21_X1 port map( B1 => n2947, B2 => n2948, A => n2809, ZN => n2946
                           );
   U2531 : NOR4_X1 port map( A1 => n2949, A2 => n2950, A3 => n2951, A4 => n2952
                           , ZN => n2948);
   U2532 : OAI221_X1 port map( B1 => n2141, B2 => n2814, C1 => n2253, C2 => 
                           n2815, A => n2953, ZN => n2952);
   U2533 : AOI22_X1 port map( A1 => n2817, A2 => n3406, B1 => n2818, B2 => 
                           n3414, ZN => n2953);
   U2534 : OAI221_X1 port map( B1 => n2142, B2 => n2819, C1 => n2261, C2 => 
                           n2820, A => n2954, ZN => n2951);
   U2535 : AOI22_X1 port map( A1 => n2822, A2 => n3470, B1 => n2823, B2 => 
                           n3478, ZN => n2954);
   U2536 : OAI221_X1 port map( B1 => n2117, B2 => n2824, C1 => n2208, C2 => 
                           n2825, A => n2955, ZN => n2950);
   U2537 : AOI22_X1 port map( A1 => n2827, A2 => n2088, B1 => n2828, B2 => 
                           n2195, ZN => n2955);
   U2538 : OAI221_X1 port map( B1 => n2118, B2 => n2829, C1 => n2209, C2 => 
                           n2830, A => n2956, ZN => n2949);
   U2539 : AOI22_X1 port map( A1 => n2832, A2 => n3374, B1 => n2833, B2 => 
                           n3382, ZN => n2956);
   U2540 : NOR4_X1 port map( A1 => n2957, A2 => n2958, A3 => n2959, A4 => n2960
                           , ZN => n2947);
   U2541 : OAI221_X1 port map( B1 => n2128, B2 => n2838, C1 => n2277, C2 => 
                           n2839, A => n2961, ZN => n2960);
   U2542 : AOI22_X1 port map( A1 => n2841, A2 => n3430, B1 => n2842, B2 => 
                           n3422, ZN => n2961);
   U2543 : OAI221_X1 port map( B1 => n2152, B2 => n2843, C1 => n2269, C2 => 
                           n2844, A => n2962, ZN => n2959);
   U2544 : AOI22_X1 port map( A1 => n2846, A2 => n3494, B1 => n2847, B2 => 
                           n3486, ZN => n2962);
   U2545 : OAI221_X1 port map( B1 => n2096, B2 => n2848, C1 => n2228, C2 => 
                           n2849, A => n2963, ZN => n2958);
   U2546 : AOI22_X1 port map( A1 => n2851, A2 => n3286, B1 => n2852, B2 => 
                           n3278, ZN => n2963);
   U2547 : OAI221_X1 port map( B1 => n2104, B2 => n2853, C1 => n2219, C2 => 
                           n2854, A => n2964, ZN => n2957);
   U2548 : AOI22_X1 port map( A1 => n2856, A2 => n3334, B1 => n2857, B2 => 
                           n3326, ZN => n2964);
   U2549 : AOI22_X1 port map( A1 => n2858, A2 => n3518, B1 => n2859, B2 => 
                           n2245, ZN => n2944);
   U2550 : OAI21_X1 port map( B1 => n2801, B2 => n2341, A => n2374, ZN => n1447
                           );
   U2551 : OAI211_X1 port map( C1 => n2801, C2 => n2366, A => n2965, B => n2966
                           , ZN => n1446);
   U2552 : AOI221_X1 port map( B1 => n2804, B2 => n3528, C1 => n2805, C2 => 
                           n2237, A => n2967, ZN => n2966);
   U2553 : AOI21_X1 port map( B1 => n2968, B2 => n2969, A => n2809, ZN => n2967
                           );
   U2554 : NOR4_X1 port map( A1 => n2970, A2 => n2971, A3 => n2972, A4 => n2973
                           , ZN => n2969);
   U2555 : OAI221_X1 port map( B1 => n2143, B2 => n2814, C1 => n2254, C2 => 
                           n2815, A => n2974, ZN => n2973);
   U2556 : AOI22_X1 port map( A1 => n2817, A2 => n3408, B1 => n2818, B2 => 
                           n3416, ZN => n2974);
   U2557 : OAI221_X1 port map( B1 => n2144, B2 => n2819, C1 => n2262, C2 => 
                           n2820, A => n2975, ZN => n2972);
   U2558 : AOI22_X1 port map( A1 => n2822, A2 => n3472, B1 => n2823, B2 => 
                           n3480, ZN => n2975);
   U2559 : OAI221_X1 port map( B1 => n2119, B2 => n2824, C1 => n2210, C2 => 
                           n2825, A => n2976, ZN => n2971);
   U2560 : AOI22_X1 port map( A1 => n2827, A2 => n2089, B1 => n2828, B2 => 
                           n2196, ZN => n2976);
   U2561 : OAI221_X1 port map( B1 => n2120, B2 => n2829, C1 => n2211, C2 => 
                           n2830, A => n2977, ZN => n2970);
   U2562 : AOI22_X1 port map( A1 => n2832, A2 => n3376, B1 => n2833, B2 => 
                           n3384, ZN => n2977);
   U2563 : NOR4_X1 port map( A1 => n2978, A2 => n2979, A3 => n2980, A4 => n2981
                           , ZN => n2968);
   U2564 : OAI221_X1 port map( B1 => n2129, B2 => n2838, C1 => n2278, C2 => 
                           n2839, A => n2982, ZN => n2981);
   U2565 : AOI22_X1 port map( A1 => n2841, A2 => n3432, B1 => n2842, B2 => 
                           n3424, ZN => n2982);
   U2566 : OAI221_X1 port map( B1 => n2153, B2 => n2843, C1 => n2270, C2 => 
                           n2844, A => n2983, ZN => n2980);
   U2567 : AOI22_X1 port map( A1 => n2846, A2 => n3496, B1 => n2847, B2 => 
                           n3488, ZN => n2983);
   U2568 : OAI221_X1 port map( B1 => n2097, B2 => n2848, C1 => n2229, C2 => 
                           n2849, A => n2984, ZN => n2979);
   U2569 : AOI22_X1 port map( A1 => n2851, A2 => n3288, B1 => n2852, B2 => 
                           n3280, ZN => n2984);
   U2570 : OAI221_X1 port map( B1 => n2105, B2 => n2853, C1 => n2220, C2 => 
                           n2854, A => n2985, ZN => n2978);
   U2571 : AOI22_X1 port map( A1 => n2856, A2 => n3336, B1 => n2857, B2 => 
                           n3328, ZN => n2985);
   U2572 : AOI22_X1 port map( A1 => n2858, A2 => n3520, B1 => n2859, B2 => 
                           n2246, ZN => n2965);
   U2573 : OAI21_X1 port map( B1 => n2801, B2 => n2342, A => n2374, ZN => n1445
                           );
   U2574 : OAI211_X1 port map( C1 => n2801, C2 => n2367, A => n2986, B => n2987
                           , ZN => n1444);
   U2575 : AOI221_X1 port map( B1 => n2804, B2 => n3527, C1 => n2805, C2 => 
                           n2238, A => n2988, ZN => n2987);
   U2576 : AOI21_X1 port map( B1 => n2989, B2 => n2990, A => n2809, ZN => n2988
                           );
   U2577 : OAI21_X1 port map( B1 => n2991, B2 => n2992, A => n2801, ZN => n2809
                           );
   U2578 : NOR4_X1 port map( A1 => n2993, A2 => n2994, A3 => n2995, A4 => n2996
                           , ZN => n2990);
   U2579 : OAI221_X1 port map( B1 => n2145, B2 => n2814, C1 => n2255, C2 => 
                           n2815, A => n2997, ZN => n2996);
   U2580 : AOI22_X1 port map( A1 => n2817, A2 => n3407, B1 => n2818, B2 => 
                           n3415, ZN => n2997);
   U2581 : AND2_X1 port map( A1 => n2998, A2 => n2999, ZN => n2818);
   U2582 : AND2_X1 port map( A1 => n3000, A2 => n2999, ZN => n2817);
   U2583 : NAND2_X1 port map( A1 => n2998, A2 => n3001, ZN => n2815);
   U2584 : NAND2_X1 port map( A1 => n3000, A2 => n3001, ZN => n2814);
   U2585 : OAI221_X1 port map( B1 => n2146, B2 => n2819, C1 => n2263, C2 => 
                           n2820, A => n3002, ZN => n2995);
   U2586 : AOI22_X1 port map( A1 => n2822, A2 => n3471, B1 => n2823, B2 => 
                           n3479, ZN => n3002);
   U2587 : AND2_X1 port map( A1 => n3003, A2 => n2999, ZN => n2823);
   U2588 : AND2_X1 port map( A1 => n3004, A2 => n2999, ZN => n2822);
   U2589 : NAND2_X1 port map( A1 => n3003, A2 => n3001, ZN => n2820);
   U2590 : NAND2_X1 port map( A1 => n3004, A2 => n3001, ZN => n2819);
   U2591 : OAI221_X1 port map( B1 => n2121, B2 => n2824, C1 => n2212, C2 => 
                           n2825, A => n3005, ZN => n2994);
   U2592 : AOI22_X1 port map( A1 => n2827, A2 => n2090, B1 => n2828, B2 => 
                           n2197, ZN => n3005);
   U2593 : AND2_X1 port map( A1 => n3006, A2 => n3007, ZN => n2828);
   U2594 : AND2_X1 port map( A1 => n3006, A2 => n3008, ZN => n2827);
   U2595 : NAND2_X1 port map( A1 => n3007, A2 => n3001, ZN => n2825);
   U2596 : NAND2_X1 port map( A1 => n3008, A2 => n3001, ZN => n2824);
   U2597 : OAI221_X1 port map( B1 => n2122, B2 => n2829, C1 => n2213, C2 => 
                           n2830, A => n3009, ZN => n2993);
   U2598 : AOI22_X1 port map( A1 => n2832, A2 => n3375, B1 => n2833, B2 => 
                           n3383, ZN => n3009);
   U2599 : AND2_X1 port map( A1 => n3001, A2 => n3010, ZN => n2833);
   U2600 : AND2_X1 port map( A1 => n3001, A2 => n3011, ZN => n2832);
   U2601 : NOR2_X1 port map( A1 => N1726, A2 => N1727, ZN => n3001);
   U2602 : NAND2_X1 port map( A1 => n3010, A2 => n2999, ZN => n2830);
   U2603 : NAND2_X1 port map( A1 => n2999, A2 => n3011, ZN => n2829);
   U2604 : NOR4_X1 port map( A1 => n3012, A2 => n3013, A3 => n3014, A4 => n3015
                           , ZN => n2989);
   U2605 : OAI221_X1 port map( B1 => n2130, B2 => n2838, C1 => n2279, C2 => 
                           n2839, A => n3016, ZN => n3015);
   U2606 : AOI22_X1 port map( A1 => n2841, A2 => n3431, B1 => n2842, B2 => 
                           n3423, ZN => n3016);
   U2607 : AND2_X1 port map( A1 => n3017, A2 => n3000, ZN => n2842);
   U2608 : AND2_X1 port map( A1 => n3017, A2 => n2998, ZN => n2841);
   U2609 : NAND2_X1 port map( A1 => n3000, A2 => n3006, ZN => n2839);
   U2610 : NOR3_X1 port map( A1 => n2383, A2 => N1729, A3 => n2391, ZN => n3000
                           );
   U2611 : NAND2_X1 port map( A1 => n2998, A2 => n3006, ZN => n2838);
   U2612 : NOR3_X1 port map( A1 => N1725, A2 => N1729, A3 => n2391, ZN => n2998
                           );
   U2613 : OAI221_X1 port map( B1 => n2154, B2 => n2843, C1 => n2271, C2 => 
                           n2844, A => n3018, ZN => n3014);
   U2614 : AOI22_X1 port map( A1 => n2846, A2 => n3495, B1 => n2847, B2 => 
                           n3487, ZN => n3018);
   U2615 : AND2_X1 port map( A1 => n3017, A2 => n3004, ZN => n2847);
   U2616 : AND2_X1 port map( A1 => n3017, A2 => n3003, ZN => n2846);
   U2617 : NAND2_X1 port map( A1 => n3004, A2 => n3006, ZN => n2844);
   U2618 : NOR3_X1 port map( A1 => N1728, A2 => N1729, A3 => n2383, ZN => n3004
                           );
   U2619 : NAND2_X1 port map( A1 => n3003, A2 => n3006, ZN => n2843);
   U2620 : NOR3_X1 port map( A1 => N1728, A2 => N1729, A3 => N1725, ZN => n3003
                           );
   U2621 : OAI221_X1 port map( B1 => n2098, B2 => n2848, C1 => n2230, C2 => 
                           n2849, A => n3019, ZN => n3013);
   U2622 : AOI22_X1 port map( A1 => n2851, A2 => n3287, B1 => n2852, B2 => 
                           n3279, ZN => n3019);
   U2623 : AND2_X1 port map( A1 => n3008, A2 => n2999, ZN => n2852);
   U2624 : AND2_X1 port map( A1 => n3007, A2 => n2999, ZN => n2851);
   U2625 : NOR2_X1 port map( A1 => n2385, A2 => N1726, ZN => n2999);
   U2626 : NAND2_X1 port map( A1 => n3017, A2 => n3008, ZN => n2849);
   U2627 : NOR3_X1 port map( A1 => n2383, A2 => n2380, A3 => n2391, ZN => n3008
                           );
   U2628 : NAND2_X1 port map( A1 => n3017, A2 => n3007, ZN => n2848);
   U2629 : NOR3_X1 port map( A1 => n2380, A2 => N1725, A3 => n2391, ZN => n3007
                           );
   U2630 : INV_X1 port map( A => N1728, ZN => n2391);
   U2631 : OAI221_X1 port map( B1 => n2106, B2 => n2853, C1 => n2221, C2 => 
                           n2854, A => n3020, ZN => n3012);
   U2632 : AOI22_X1 port map( A1 => n2856, A2 => n3335, B1 => n2857, B2 => 
                           n3327, ZN => n3020);
   U2633 : AND2_X1 port map( A1 => n3006, A2 => n3011, ZN => n2857);
   U2634 : AND2_X1 port map( A1 => n3006, A2 => n3010, ZN => n2856);
   U2635 : NOR2_X1 port map( A1 => n2385, A2 => n2384, ZN => n3006);
   U2636 : INV_X1 port map( A => N1727, ZN => n2385);
   U2637 : NAND2_X1 port map( A1 => n3017, A2 => n3011, ZN => n2854);
   U2638 : NOR3_X1 port map( A1 => n2380, A2 => N1728, A3 => n2383, ZN => n3011
                           );
   U2639 : INV_X1 port map( A => N1725, ZN => n2383);
   U2640 : NAND2_X1 port map( A1 => n3017, A2 => n3010, ZN => n2853);
   U2641 : NOR3_X1 port map( A1 => N1725, A2 => N1728, A3 => n2380, ZN => n3010
                           );
   U2642 : INV_X1 port map( A => N1729, ZN => n2380);
   U2643 : NOR2_X1 port map( A1 => n2384, A2 => N1727, ZN => n3017);
   U2644 : INV_X1 port map( A => N1726, ZN => n2384);
   U2645 : AND3_X1 port map( A1 => n3021, A2 => n3022, A3 => n3023, ZN => n2805
                           );
   U2646 : AND3_X1 port map( A1 => n3023, A2 => n3021, A3 => ADD_RD2(1), ZN => 
                           n2804);
   U2647 : AOI22_X1 port map( A1 => n2858, A2 => n3519, B1 => n2859, B2 => 
                           n2247, ZN => n2986);
   U2648 : AND3_X1 port map( A1 => n3023, A2 => n3022, A3 => ADD_RD2(0), ZN => 
                           n2859);
   U2649 : AND3_X1 port map( A1 => ADD_RD2(1), A2 => n3023, A3 => ADD_RD2(0), 
                           ZN => n2858);
   U2650 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => n2801, A3 => ADD_RD2(3), 
                           ZN => n3023);
   U2651 : OAI21_X1 port map( B1 => n2801, B2 => n2343, A => n2374, ZN => n1443
                           );
   U2652 : NAND2_X1 port map( A1 => n3024, A2 => n2374, ZN => n2801);
   U2653 : NAND2_X1 port map( A1 => RD2, A2 => n2432, ZN => n3024);
   U2654 : NOR2_X1 port map( A1 => n3025, A2 => n2390, ZN => n2432);
   U2655 : NAND3_X1 port map( A1 => n3026, A2 => n3027, A3 => n3028, ZN => 
                           n1442);
   U2656 : AOI211_X1 port map( C1 => n3029, C2 => n3515, A => n3030, B => n3031
                           , ZN => n3028);
   U2657 : MUX2_X1 port map( A => n3032, B => n1361, S => n2471, Z => n3031);
   U2658 : NAND4_X1 port map( A1 => n3033, A2 => n3034, A3 => n3035, A4 => 
                           n3036, ZN => n3032);
   U2659 : AOI221_X1 port map( B1 => n3339, B2 => n3037, C1 => n3331, C2 => 
                           n3038, A => n3039, ZN => n3036);
   U2660 : OAI22_X1 port map( A1 => n2535, A2 => n2099, B1 => n2538, B2 => 
                           n2214, ZN => n3039);
   U2661 : AOI221_X1 port map( B1 => n3040, B2 => n2083, C1 => n3041, C2 => 
                           n2190, A => n3042, ZN => n3035);
   U2662 : OAI22_X1 port map( A1 => n2554, A2 => n2223, B1 => n2552, B2 => 
                           n2091, ZN => n3042);
   U2663 : AOI221_X1 port map( B1 => n3467, B2 => n3043, C1 => n3459, C2 => 
                           n3044, A => n3045, ZN => n3034);
   U2664 : OAI22_X1 port map( A1 => n2493, A2 => n2288, B1 => n2496, B2 => 
                           n2179, ZN => n3045);
   U2665 : AOI221_X1 port map( B1 => n3395, B2 => n3046, C1 => n3403, C2 => 
                           n3047, A => n3048, ZN => n3033);
   U2666 : OAI22_X1 port map( A1 => n2514, A2 => n2296, B1 => n2512, B2 => 
                           n2171, ZN => n3048);
   U2667 : OAI22_X1 port map( A1 => n2280, A2 => n3049, B1 => n2155, B2 => 
                           n3050, ZN => n3030);
   U2668 : AOI22_X1 port map( A1 => n3051, A2 => n3052, B1 => n3053, B2 => 
                           n3054, ZN => n3027);
   U2669 : OAI221_X1 port map( B1 => n2198, B2 => n3055, C1 => n2107, C2 => 
                           n3056, A => n3057, ZN => n3054);
   U2670 : AOI22_X1 port map( A1 => n3058, A2 => n3451, B1 => n3059, B2 => 
                           n3443, ZN => n3057);
   U2671 : OAI221_X1 port map( B1 => n2199, B2 => n3055, C1 => n2108, C2 => 
                           n3056, A => n3060, ZN => n3052);
   U2672 : AOI22_X1 port map( A1 => n3058, A2 => n3483, B1 => n3059, B2 => 
                           n3475, ZN => n3060);
   U2673 : AOI22_X1 port map( A1 => n3061, A2 => n3062, B1 => n3063, B2 => 
                           n3507, ZN => n3026);
   U2674 : OAI221_X1 port map( B1 => n2163, B2 => n3055, C1 => n2304, C2 => 
                           n3056, A => n3064, ZN => n3062);
   U2675 : AOI22_X1 port map( A1 => n3058, A2 => n3419, B1 => n3059, B2 => 
                           n3411, ZN => n3064);
   U2676 : OAI21_X1 port map( B1 => n3065, B2 => n2344, A => n3066, ZN => n1441
                           );
   U2677 : NAND3_X1 port map( A1 => n3067, A2 => n3068, A3 => n3069, ZN => 
                           n1440);
   U2678 : AOI211_X1 port map( C1 => n3029, C2 => n3508, A => n3070, B => n3071
                           , ZN => n3069);
   U2679 : MUX2_X1 port map( A => n3072, B => n1363, S => n2471, Z => n3071);
   U2680 : NAND4_X1 port map( A1 => n3073, A2 => n3074, A3 => n3075, A4 => 
                           n3076, ZN => n3072);
   U2681 : AOI221_X1 port map( B1 => n3332, B2 => n3037, C1 => n3324, C2 => 
                           n3038, A => n3077, ZN => n3076);
   U2682 : OAI22_X1 port map( A1 => n2535, A2 => n2100, B1 => n2538, B2 => 
                           n2215, ZN => n3077);
   U2683 : AOI221_X1 port map( B1 => n3040, B2 => n2084, C1 => n3041, C2 => 
                           n2191, A => n3078, ZN => n3075);
   U2684 : OAI22_X1 port map( A1 => n2554, A2 => n2224, B1 => n2552, B2 => 
                           n2092, ZN => n3078);
   U2685 : AOI221_X1 port map( B1 => n3460, B2 => n3043, C1 => n3452, C2 => 
                           n3044, A => n3079, ZN => n3074);
   U2686 : OAI22_X1 port map( A1 => n2493, A2 => n2289, B1 => n2496, B2 => 
                           n2180, ZN => n3079);
   U2687 : AOI221_X1 port map( B1 => n3388, B2 => n3046, C1 => n3396, C2 => 
                           n3047, A => n3080, ZN => n3073);
   U2688 : OAI22_X1 port map( A1 => n2514, A2 => n2297, B1 => n2512, B2 => 
                           n2172, ZN => n3080);
   U2689 : OAI22_X1 port map( A1 => n2281, A2 => n3049, B1 => n2156, B2 => 
                           n3050, ZN => n3070);
   U2690 : AOI22_X1 port map( A1 => n3051, A2 => n3081, B1 => n3053, B2 => 
                           n3082, ZN => n3068);
   U2691 : OAI221_X1 port map( B1 => n2200, B2 => n3055, C1 => n2109, C2 => 
                           n3056, A => n3083, ZN => n3082);
   U2692 : AOI22_X1 port map( A1 => n3058, A2 => n3444, B1 => n3059, B2 => 
                           n3436, ZN => n3083);
   U2693 : OAI221_X1 port map( B1 => n2201, B2 => n3055, C1 => n2110, C2 => 
                           n3056, A => n3084, ZN => n3081);
   U2694 : AOI22_X1 port map( A1 => n3058, A2 => n3476, B1 => n3059, B2 => 
                           n3468, ZN => n3084);
   U2695 : AOI22_X1 port map( A1 => n3061, A2 => n3085, B1 => n3063, B2 => 
                           n3500, ZN => n3067);
   U2696 : OAI221_X1 port map( B1 => n2164, B2 => n3055, C1 => n2305, C2 => 
                           n3056, A => n3086, ZN => n3085);
   U2697 : AOI22_X1 port map( A1 => n3058, A2 => n3412, B1 => n3059, B2 => 
                           n3404, ZN => n3086);
   U2698 : OAI21_X1 port map( B1 => n3065, B2 => n2345, A => n3066, ZN => n1439
                           );
   U2699 : NAND3_X1 port map( A1 => n3087, A2 => n3088, A3 => n3089, ZN => 
                           n1438);
   U2700 : AOI211_X1 port map( C1 => n3029, C2 => n3514, A => n3090, B => n3091
                           , ZN => n3089);
   U2701 : MUX2_X1 port map( A => n3092, B => n1365, S => n2471, Z => n3091);
   U2702 : NAND4_X1 port map( A1 => n3093, A2 => n3094, A3 => n3095, A4 => 
                           n3096, ZN => n3092);
   U2703 : AOI221_X1 port map( B1 => n3338, B2 => n3037, C1 => n3330, C2 => 
                           n3038, A => n3097, ZN => n3096);
   U2704 : OAI22_X1 port map( A1 => n2535, A2 => n2101, B1 => n2538, B2 => 
                           n2216, ZN => n3097);
   U2705 : AOI221_X1 port map( B1 => n3040, B2 => n2085, C1 => n3041, C2 => 
                           n2192, A => n3098, ZN => n3095);
   U2706 : OAI22_X1 port map( A1 => n2554, A2 => n2225, B1 => n2552, B2 => 
                           n2093, ZN => n3098);
   U2707 : AOI221_X1 port map( B1 => n3466, B2 => n3043, C1 => n3458, C2 => 
                           n3044, A => n3099, ZN => n3094);
   U2708 : OAI22_X1 port map( A1 => n2493, A2 => n2290, B1 => n2496, B2 => 
                           n2181, ZN => n3099);
   U2709 : AOI221_X1 port map( B1 => n3394, B2 => n3046, C1 => n3402, C2 => 
                           n3047, A => n3100, ZN => n3093);
   U2710 : OAI22_X1 port map( A1 => n2514, A2 => n2298, B1 => n2512, B2 => 
                           n2173, ZN => n3100);
   U2711 : OAI22_X1 port map( A1 => n2282, A2 => n3049, B1 => n2157, B2 => 
                           n3050, ZN => n3090);
   U2712 : AOI22_X1 port map( A1 => n3051, A2 => n3101, B1 => n3053, B2 => 
                           n3102, ZN => n3088);
   U2713 : OAI221_X1 port map( B1 => n2202, B2 => n3055, C1 => n2111, C2 => 
                           n3056, A => n3103, ZN => n3102);
   U2714 : AOI22_X1 port map( A1 => n3058, A2 => n3450, B1 => n3059, B2 => 
                           n3442, ZN => n3103);
   U2715 : OAI221_X1 port map( B1 => n2203, B2 => n3055, C1 => n2112, C2 => 
                           n3056, A => n3104, ZN => n3101);
   U2716 : AOI22_X1 port map( A1 => n3058, A2 => n3482, B1 => n3059, B2 => 
                           n3474, ZN => n3104);
   U2717 : AOI22_X1 port map( A1 => n3061, A2 => n3105, B1 => n3063, B2 => 
                           n3506, ZN => n3087);
   U2718 : OAI221_X1 port map( B1 => n2165, B2 => n3055, C1 => n2306, C2 => 
                           n3056, A => n3106, ZN => n3105);
   U2719 : AOI22_X1 port map( A1 => n3058, A2 => n3418, B1 => n3059, B2 => 
                           n3410, ZN => n3106);
   U2720 : OAI21_X1 port map( B1 => n3065, B2 => n2346, A => n3066, ZN => n1437
                           );
   U2721 : NAND3_X1 port map( A1 => n3107, A2 => n3108, A3 => n3109, ZN => 
                           n1436);
   U2722 : AOI211_X1 port map( C1 => n3029, C2 => n3509, A => n3110, B => n3111
                           , ZN => n3109);
   U2723 : MUX2_X1 port map( A => n3112, B => n1367, S => n2471, Z => n3111);
   U2724 : NAND4_X1 port map( A1 => n3113, A2 => n3114, A3 => n3115, A4 => 
                           n3116, ZN => n3112);
   U2725 : AOI221_X1 port map( B1 => n3333, B2 => n3037, C1 => n3325, C2 => 
                           n3038, A => n3117, ZN => n3116);
   U2726 : OAI22_X1 port map( A1 => n2535, A2 => n2102, B1 => n2538, B2 => 
                           n2217, ZN => n3117);
   U2727 : AOI221_X1 port map( B1 => n3040, B2 => n2086, C1 => n3041, C2 => 
                           n2193, A => n3118, ZN => n3115);
   U2728 : OAI22_X1 port map( A1 => n2554, A2 => n2226, B1 => n2552, B2 => 
                           n2094, ZN => n3118);
   U2729 : AOI221_X1 port map( B1 => n3461, B2 => n3043, C1 => n3453, C2 => 
                           n3044, A => n3119, ZN => n3114);
   U2730 : OAI22_X1 port map( A1 => n2493, A2 => n2291, B1 => n2496, B2 => 
                           n2182, ZN => n3119);
   U2731 : AOI221_X1 port map( B1 => n3389, B2 => n3046, C1 => n3397, C2 => 
                           n3047, A => n3120, ZN => n3113);
   U2732 : OAI22_X1 port map( A1 => n2514, A2 => n2299, B1 => n2512, B2 => 
                           n2174, ZN => n3120);
   U2733 : OAI22_X1 port map( A1 => n2283, A2 => n3049, B1 => n2158, B2 => 
                           n3050, ZN => n3110);
   U2734 : AOI22_X1 port map( A1 => n3051, A2 => n3121, B1 => n3053, B2 => 
                           n3122, ZN => n3108);
   U2735 : OAI221_X1 port map( B1 => n2204, B2 => n3055, C1 => n2113, C2 => 
                           n3056, A => n3123, ZN => n3122);
   U2736 : AOI22_X1 port map( A1 => n3058, A2 => n3445, B1 => n3059, B2 => 
                           n3437, ZN => n3123);
   U2737 : OAI221_X1 port map( B1 => n2205, B2 => n3055, C1 => n2114, C2 => 
                           n3056, A => n3124, ZN => n3121);
   U2738 : AOI22_X1 port map( A1 => n3058, A2 => n3477, B1 => n3059, B2 => 
                           n3469, ZN => n3124);
   U2739 : AOI22_X1 port map( A1 => n3061, A2 => n3125, B1 => n3063, B2 => 
                           n3501, ZN => n3107);
   U2740 : OAI221_X1 port map( B1 => n2166, B2 => n3055, C1 => n2307, C2 => 
                           n3056, A => n3126, ZN => n3125);
   U2741 : AOI22_X1 port map( A1 => n3058, A2 => n3413, B1 => n3059, B2 => 
                           n3405, ZN => n3126);
   U2742 : OAI21_X1 port map( B1 => n3065, B2 => n2347, A => n3066, ZN => n1435
                           );
   U2743 : NAND3_X1 port map( A1 => n3127, A2 => n3128, A3 => n3129, ZN => 
                           n1434);
   U2744 : AOI211_X1 port map( C1 => n3029, C2 => n3513, A => n3130, B => n3131
                           , ZN => n3129);
   U2745 : MUX2_X1 port map( A => n3132, B => n1369, S => n2471, Z => n3131);
   U2746 : NAND4_X1 port map( A1 => n3133, A2 => n3134, A3 => n3135, A4 => 
                           n3136, ZN => n3132);
   U2747 : AOI221_X1 port map( B1 => n3337, B2 => n3037, C1 => n3329, C2 => 
                           n3038, A => n3137, ZN => n3136);
   U2748 : OAI22_X1 port map( A1 => n2535, A2 => n2103, B1 => n2538, B2 => 
                           n2218, ZN => n3137);
   U2749 : AOI221_X1 port map( B1 => n3040, B2 => n2087, C1 => n3041, C2 => 
                           n2194, A => n3138, ZN => n3135);
   U2750 : OAI22_X1 port map( A1 => n2554, A2 => n2227, B1 => n2552, B2 => 
                           n2095, ZN => n3138);
   U2751 : AOI221_X1 port map( B1 => n3465, B2 => n3043, C1 => n3457, C2 => 
                           n3044, A => n3139, ZN => n3134);
   U2752 : OAI22_X1 port map( A1 => n2493, A2 => n2292, B1 => n2496, B2 => 
                           n2183, ZN => n3139);
   U2753 : AOI221_X1 port map( B1 => n3393, B2 => n3046, C1 => n3401, C2 => 
                           n3047, A => n3140, ZN => n3133);
   U2754 : OAI22_X1 port map( A1 => n2514, A2 => n2300, B1 => n2512, B2 => 
                           n2175, ZN => n3140);
   U2755 : OAI22_X1 port map( A1 => n2284, A2 => n3049, B1 => n2159, B2 => 
                           n3050, ZN => n3130);
   U2756 : AOI22_X1 port map( A1 => n3051, A2 => n3141, B1 => n3053, B2 => 
                           n3142, ZN => n3128);
   U2757 : OAI221_X1 port map( B1 => n2206, B2 => n3055, C1 => n2115, C2 => 
                           n3056, A => n3143, ZN => n3142);
   U2758 : AOI22_X1 port map( A1 => n3058, A2 => n3449, B1 => n3059, B2 => 
                           n3441, ZN => n3143);
   U2759 : OAI221_X1 port map( B1 => n2207, B2 => n3055, C1 => n2116, C2 => 
                           n3056, A => n3144, ZN => n3141);
   U2760 : AOI22_X1 port map( A1 => n3058, A2 => n3481, B1 => n3059, B2 => 
                           n3473, ZN => n3144);
   U2761 : AOI22_X1 port map( A1 => n3061, A2 => n3145, B1 => n3063, B2 => 
                           n3505, ZN => n3127);
   U2762 : OAI221_X1 port map( B1 => n2167, B2 => n3055, C1 => n2308, C2 => 
                           n3056, A => n3146, ZN => n3145);
   U2763 : AOI22_X1 port map( A1 => n3058, A2 => n3417, B1 => n3059, B2 => 
                           n3409, ZN => n3146);
   U2764 : OAI21_X1 port map( B1 => n3065, B2 => n2348, A => n3066, ZN => n1433
                           );
   U2765 : NAND3_X1 port map( A1 => n3147, A2 => n3148, A3 => n3149, ZN => 
                           n1432);
   U2766 : AOI211_X1 port map( C1 => n3029, C2 => n3510, A => n3150, B => n3151
                           , ZN => n3149);
   U2767 : MUX2_X1 port map( A => n3152, B => n1371, S => n2471, Z => n3151);
   U2768 : NAND4_X1 port map( A1 => n3153, A2 => n3154, A3 => n3155, A4 => 
                           n3156, ZN => n3152);
   U2769 : AOI221_X1 port map( B1 => n3334, B2 => n3037, C1 => n3326, C2 => 
                           n3038, A => n3157, ZN => n3156);
   U2770 : OAI22_X1 port map( A1 => n2535, A2 => n2104, B1 => n2538, B2 => 
                           n2219, ZN => n3157);
   U2771 : AOI221_X1 port map( B1 => n3040, B2 => n2088, C1 => n3041, C2 => 
                           n2195, A => n3158, ZN => n3155);
   U2772 : OAI22_X1 port map( A1 => n2554, A2 => n2228, B1 => n2552, B2 => 
                           n2096, ZN => n3158);
   U2773 : AOI221_X1 port map( B1 => n3462, B2 => n3043, C1 => n3454, C2 => 
                           n3044, A => n3159, ZN => n3154);
   U2774 : OAI22_X1 port map( A1 => n2493, A2 => n2293, B1 => n2496, B2 => 
                           n2184, ZN => n3159);
   U2775 : AOI221_X1 port map( B1 => n3390, B2 => n3046, C1 => n3398, C2 => 
                           n3047, A => n3160, ZN => n3153);
   U2776 : OAI22_X1 port map( A1 => n2514, A2 => n2301, B1 => n2512, B2 => 
                           n2176, ZN => n3160);
   U2777 : OAI22_X1 port map( A1 => n2285, A2 => n3049, B1 => n2160, B2 => 
                           n3050, ZN => n3150);
   U2778 : AOI22_X1 port map( A1 => n3051, A2 => n3161, B1 => n3053, B2 => 
                           n3162, ZN => n3148);
   U2779 : OAI221_X1 port map( B1 => n2208, B2 => n3055, C1 => n2117, C2 => 
                           n3056, A => n3163, ZN => n3162);
   U2780 : AOI22_X1 port map( A1 => n3058, A2 => n3446, B1 => n3059, B2 => 
                           n3438, ZN => n3163);
   U2781 : OAI221_X1 port map( B1 => n2209, B2 => n3055, C1 => n2118, C2 => 
                           n3056, A => n3164, ZN => n3161);
   U2782 : AOI22_X1 port map( A1 => n3058, A2 => n3478, B1 => n3059, B2 => 
                           n3470, ZN => n3164);
   U2783 : AOI22_X1 port map( A1 => n3061, A2 => n3165, B1 => n3063, B2 => 
                           n3502, ZN => n3147);
   U2784 : OAI221_X1 port map( B1 => n2168, B2 => n3055, C1 => n2309, C2 => 
                           n3056, A => n3166, ZN => n3165);
   U2785 : AOI22_X1 port map( A1 => n3058, A2 => n3414, B1 => n3059, B2 => 
                           n3406, ZN => n3166);
   U2786 : OAI21_X1 port map( B1 => n3065, B2 => n2349, A => n3066, ZN => n1431
                           );
   U2787 : NAND3_X1 port map( A1 => n3167, A2 => n3168, A3 => n3169, ZN => 
                           n1430);
   U2788 : AOI211_X1 port map( C1 => n3029, C2 => n3512, A => n3170, B => n3171
                           , ZN => n3169);
   U2789 : MUX2_X1 port map( A => n3172, B => n1373, S => n2471, Z => n3171);
   U2790 : NAND4_X1 port map( A1 => n3173, A2 => n3174, A3 => n3175, A4 => 
                           n3176, ZN => n3172);
   U2791 : AOI221_X1 port map( B1 => n3336, B2 => n3037, C1 => n3328, C2 => 
                           n3038, A => n3177, ZN => n3176);
   U2792 : OAI22_X1 port map( A1 => n2535, A2 => n2105, B1 => n2538, B2 => 
                           n2220, ZN => n3177);
   U2793 : AOI221_X1 port map( B1 => n3040, B2 => n2089, C1 => n3041, C2 => 
                           n2196, A => n3178, ZN => n3175);
   U2794 : OAI22_X1 port map( A1 => n2554, A2 => n2229, B1 => n2552, B2 => 
                           n2097, ZN => n3178);
   U2795 : AOI221_X1 port map( B1 => n3464, B2 => n3043, C1 => n3456, C2 => 
                           n3044, A => n3179, ZN => n3174);
   U2796 : OAI22_X1 port map( A1 => n2493, A2 => n2294, B1 => n2496, B2 => 
                           n2185, ZN => n3179);
   U2797 : AOI221_X1 port map( B1 => n3392, B2 => n3046, C1 => n3400, C2 => 
                           n3047, A => n3180, ZN => n3173);
   U2798 : OAI22_X1 port map( A1 => n2514, A2 => n2302, B1 => n2512, B2 => 
                           n2177, ZN => n3180);
   U2799 : OAI22_X1 port map( A1 => n2286, A2 => n3049, B1 => n2161, B2 => 
                           n3050, ZN => n3170);
   U2800 : AOI22_X1 port map( A1 => n3051, A2 => n3181, B1 => n3053, B2 => 
                           n3182, ZN => n3168);
   U2801 : OAI221_X1 port map( B1 => n2210, B2 => n3055, C1 => n2119, C2 => 
                           n3056, A => n3183, ZN => n3182);
   U2802 : AOI22_X1 port map( A1 => n3058, A2 => n3448, B1 => n3059, B2 => 
                           n3440, ZN => n3183);
   U2803 : OAI221_X1 port map( B1 => n2211, B2 => n3055, C1 => n2120, C2 => 
                           n3056, A => n3184, ZN => n3181);
   U2804 : AOI22_X1 port map( A1 => n3058, A2 => n3480, B1 => n3059, B2 => 
                           n3472, ZN => n3184);
   U2805 : AOI22_X1 port map( A1 => n3061, A2 => n3185, B1 => n3063, B2 => 
                           n3504, ZN => n3167);
   U2806 : OAI221_X1 port map( B1 => n2169, B2 => n3055, C1 => n2310, C2 => 
                           n3056, A => n3186, ZN => n3185);
   U2807 : AOI22_X1 port map( A1 => n3058, A2 => n3416, B1 => n3059, B2 => 
                           n3408, ZN => n3186);
   U2808 : OAI21_X1 port map( B1 => n3065, B2 => n2350, A => n3066, ZN => n1429
                           );
   U2809 : NAND3_X1 port map( A1 => n3187, A2 => n3188, A3 => n3189, ZN => 
                           n1428);
   U2810 : AOI211_X1 port map( C1 => n3029, C2 => n3511, A => n3190, B => n3191
                           , ZN => n3189);
   U2811 : MUX2_X1 port map( A => n3192, B => n1375, S => n2471, Z => n3191);
   U2812 : NAND4_X1 port map( A1 => n3193, A2 => n3194, A3 => n3195, A4 => 
                           n3196, ZN => n3192);
   U2813 : AOI221_X1 port map( B1 => n3335, B2 => n3037, C1 => n3327, C2 => 
                           n3038, A => n3197, ZN => n3196);
   U2814 : OAI22_X1 port map( A1 => n2535, A2 => n2106, B1 => n2538, B2 => 
                           n2221, ZN => n3197);
   U2815 : NAND2_X1 port map( A1 => n3198, A2 => n3199, ZN => n2538);
   U2816 : NAND2_X1 port map( A1 => n3198, A2 => n3200, ZN => n2535);
   U2817 : INV_X1 port map( A => n2548, ZN => n3038);
   U2818 : NAND2_X1 port map( A1 => n3201, A2 => n3051, ZN => n2548);
   U2819 : INV_X1 port map( A => n2546, ZN => n3037);
   U2820 : NAND2_X1 port map( A1 => n3202, A2 => n3051, ZN => n2546);
   U2821 : AOI221_X1 port map( B1 => n3040, B2 => n2090, C1 => n3041, C2 => 
                           n2197, A => n3203, ZN => n3195);
   U2822 : OAI22_X1 port map( A1 => n2554, A2 => n2230, B1 => n2552, B2 => 
                           n2098, ZN => n3203);
   U2823 : NAND2_X1 port map( A1 => n3202, A2 => n3053, ZN => n2552);
   U2824 : NAND2_X1 port map( A1 => n3201, A2 => n3053, ZN => n2554);
   U2825 : INV_X1 port map( A => n2560, ZN => n3041);
   U2826 : NAND2_X1 port map( A1 => n3202, A2 => n3061, ZN => n2560);
   U2827 : AND2_X1 port map( A1 => n3200, A2 => n3585, ZN => n3202);
   U2828 : INV_X1 port map( A => n2569, ZN => n3040);
   U2829 : NAND2_X1 port map( A1 => n3201, A2 => n3061, ZN => n2569);
   U2830 : AND2_X1 port map( A1 => n3199, A2 => n3585, ZN => n3201);
   U2831 : AOI221_X1 port map( B1 => n3463, B2 => n3043, C1 => n3455, C2 => 
                           n3044, A => n3204, ZN => n3194);
   U2832 : OAI22_X1 port map( A1 => n2493, A2 => n2295, B1 => n2496, B2 => 
                           n2186, ZN => n3204);
   U2833 : NAND2_X1 port map( A1 => n3199, A2 => n3205, ZN => n2496);
   U2834 : NAND2_X1 port map( A1 => n3200, A2 => n3205, ZN => n2493);
   U2835 : INV_X1 port map( A => n2506, ZN => n3044);
   U2836 : NAND2_X1 port map( A1 => n3206, A2 => n3051, ZN => n2506);
   U2837 : INV_X1 port map( A => n2504, ZN => n3043);
   U2838 : NAND2_X1 port map( A1 => n3207, A2 => n3051, ZN => n2504);
   U2839 : AOI221_X1 port map( B1 => n3391, B2 => n3046, C1 => n3399, C2 => 
                           n3047, A => n3208, ZN => n3193);
   U2840 : OAI22_X1 port map( A1 => n2514, A2 => n2303, B1 => n2512, B2 => 
                           n2178, ZN => n3208);
   U2841 : NAND2_X1 port map( A1 => n3053, A2 => n3207, ZN => n2512);
   U2842 : NAND2_X1 port map( A1 => n3053, A2 => n3206, ZN => n2514);
   U2843 : INV_X1 port map( A => n2523, ZN => n3047);
   U2844 : NAND2_X1 port map( A1 => n3061, A2 => n3207, ZN => n2523);
   U2845 : AND2_X1 port map( A1 => n3200, A2 => n2080, ZN => n3207);
   U2846 : NOR2_X1 port map( A1 => n2082, A2 => n3589, ZN => n3200);
   U2847 : INV_X1 port map( A => n2525, ZN => n3046);
   U2848 : NAND2_X1 port map( A1 => n3061, A2 => n3206, ZN => n2525);
   U2849 : AND2_X1 port map( A1 => n3199, A2 => n2080, ZN => n3206);
   U2850 : NOR2_X1 port map( A1 => n2082, A2 => n2188, ZN => n3199);
   U2851 : OAI22_X1 port map( A1 => n2287, A2 => n3049, B1 => n2162, B2 => 
                           n3050, ZN => n3190);
   U2852 : NAND2_X1 port map( A1 => n3209, A2 => n3198, ZN => n3050);
   U2853 : NAND2_X1 port map( A1 => n3210, A2 => n3198, ZN => n3049);
   U2854 : INV_X1 port map( A => n2530, ZN => n3198);
   U2855 : NAND3_X1 port map( A1 => n2187, A2 => n2081, A3 => n3585, ZN => 
                           n2530);
   U2856 : AND2_X1 port map( A1 => n3210, A2 => n3205, ZN => n3029);
   U2857 : AOI22_X1 port map( A1 => n3051, A2 => n3211, B1 => n3053, B2 => 
                           n3212, ZN => n3188);
   U2858 : OAI221_X1 port map( B1 => n2212, B2 => n3055, C1 => n2121, C2 => 
                           n3056, A => n3213, ZN => n3212);
   U2859 : AOI22_X1 port map( A1 => n3058, A2 => n3447, B1 => n3059, B2 => 
                           n3439, ZN => n3213);
   U2860 : INV_X1 port map( A => n2508, ZN => n3053);
   U2861 : NAND2_X1 port map( A1 => n3586, A2 => n2187, ZN => n2508);
   U2862 : OAI221_X1 port map( B1 => n2213, B2 => n3055, C1 => n2122, C2 => 
                           n3056, A => n3214, ZN => n3211);
   U2863 : AOI22_X1 port map( A1 => n3058, A2 => n3479, B1 => n3059, B2 => 
                           n3471, ZN => n3214);
   U2864 : INV_X1 port map( A => n2499, ZN => n3051);
   U2865 : NAND2_X1 port map( A1 => n3587, A2 => n2081, ZN => n2499);
   U2866 : AOI22_X1 port map( A1 => n3061, A2 => n3215, B1 => n3063, B2 => 
                           n3503, ZN => n3187);
   U2867 : AND2_X1 port map( A1 => n3209, A2 => n3205, ZN => n3063);
   U2868 : INV_X1 port map( A => n2486, ZN => n3205);
   U2869 : OAI221_X1 port map( B1 => n2170, B2 => n3055, C1 => n2311, C2 => 
                           n3056, A => n3216, ZN => n3215);
   U2870 : AOI22_X1 port map( A1 => n3058, A2 => n3415, B1 => n3059, B2 => 
                           n3407, ZN => n3216);
   U2871 : AND2_X1 port map( A1 => n3209, A2 => n2080, ZN => n3059);
   U2872 : AND2_X1 port map( A1 => n3210, A2 => n2080, ZN => n3058);
   U2873 : NAND2_X1 port map( A1 => n3209, A2 => n3585, ZN => n3056);
   U2874 : NOR3_X1 port map( A1 => n2471, A2 => n3588, A3 => n2188, ZN => n3209
                           );
   U2875 : NAND2_X1 port map( A1 => n3210, A2 => n3585, ZN => n3055);
   U2876 : NOR2_X1 port map( A1 => n2557, A2 => n2471, ZN => n3210);
   U2877 : INV_X1 port map( A => n3065, ZN => n2471);
   U2878 : INV_X1 port map( A => n2516, ZN => n3061);
   U2879 : NAND2_X1 port map( A1 => n3586, A2 => n3587, ZN => n2516);
   U2880 : OAI21_X1 port map( B1 => n3065, B2 => n2351, A => n3066, ZN => n1427
                           );
   U2881 : OAI21_X1 port map( B1 => n1259, B2 => n2473, A => n2474, ZN => n1426
                           );
   U2882 : NAND3_X1 port map( A1 => n2473, A2 => n2374, A3 => n2389, ZN => 
                           n2474);
   U2883 : NAND3_X1 port map( A1 => n3217, A2 => n2374, A3 => n3218, ZN => 
                           n2473);
   U2884 : OR4_X1 port map( A1 => n2387, A2 => n2390, A3 => n2189, A4 => n3582,
                           ZN => n3218);
   U2885 : NAND4_X1 port map( A1 => n2799, A2 => n2408, A3 => n3219, A4 => 
                           n3220, ZN => n3217);
   U2886 : AOI211_X1 port map( C1 => CWP_1_port, C2 => n2082, A => n3221, B => 
                           n3222, ZN => n3220);
   U2887 : INV_X1 port map( A => n3223, ZN => n3222);
   U2888 : NAND3_X1 port map( A1 => n3224, A2 => n2399, A3 => n3225, ZN => 
                           n3221);
   U2889 : INV_X1 port map( A => n3226, ZN => n3225);
   U2890 : INV_X1 port map( A => n2407, ZN => n2399);
   U2891 : NOR3_X1 port map( A1 => n2372, A2 => n2397, A3 => n2222, ZN => n2407
                           );
   U2892 : INV_X1 port map( A => n2406, ZN => n2397);
   U2893 : NOR3_X1 port map( A1 => CWP_4_port, A2 => n2375, A3 => CWP_3_port, 
                           ZN => n2406);
   U2894 : NAND2_X1 port map( A1 => n3227, A2 => n3228, ZN => n2372);
   U2895 : NOR4_X1 port map( A1 => n3229, A2 => n3230, A3 => n3231, A4 => n3232
                           , ZN => n3228);
   U2896 : NAND4_X1 port map( A1 => n3565, A2 => n3566, A3 => n3567, A4 => 
                           n3568, ZN => n3232);
   U2897 : NAND4_X1 port map( A1 => n3569, A2 => n3570, A3 => n3571, A4 => 
                           n3572, ZN => n3231);
   U2898 : NAND4_X1 port map( A1 => n3573, A2 => n3574, A3 => n3575, A4 => 
                           n3576, ZN => n3230);
   U2899 : NAND4_X1 port map( A1 => n3577, A2 => n3578, A3 => n3579, A4 => 
                           n3580, ZN => n3229);
   U2900 : NOR4_X1 port map( A1 => n3233, A2 => n3234, A3 => n3235, A4 => n3236
                           , ZN => n3227);
   U2901 : NAND4_X1 port map( A1 => n3549, A2 => n3550, A3 => n3551, A4 => 
                           n3552, ZN => n3236);
   U2902 : NAND4_X1 port map( A1 => n3553, A2 => n3554, A3 => n3555, A4 => 
                           n3556, ZN => n3235);
   U2903 : NAND4_X1 port map( A1 => n3557, A2 => n3558, A3 => n3559, A4 => 
                           n3560, ZN => n3234);
   U2904 : NAND4_X1 port map( A1 => n3561, A2 => n3562, A3 => n3563, A4 => 
                           n3564, ZN => n3233);
   U2905 : AOI21_X1 port map( B1 => CWP_0_port, B2 => n3237, A => n3238, ZN => 
                           n3219);
   U2906 : NOR3_X1 port map( A1 => CALL, A2 => n3548, A3 => n2400, ZN => n2408)
                           ;
   U2907 : INV_X1 port map( A => n2762, ZN => n2799);
   U2908 : OAI21_X1 port map( B1 => n3239, B2 => n3240, A => n3241, ZN => n2762
                           );
   U2909 : NAND4_X1 port map( A1 => n3242, A2 => n3223, A3 => n3243, A4 => 
                           n3224, ZN => n3241);
   U2910 : NAND3_X1 port map( A1 => n3244, A2 => n2081, A3 => n3245, ZN => 
                           n3224);
   U2911 : OAI21_X1 port map( B1 => n3226, B2 => n3246, A => n3247, ZN => n3243
                           );
   U2912 : OAI22_X1 port map( A1 => n3248, A2 => n3249, B1 => n3239, B2 => 
                           n3250, ZN => n3247);
   U2913 : AOI22_X1 port map( A1 => n3251, A2 => n2081, B1 => n3245, B2 => 
                           n2187, ZN => n3250);
   U2914 : NAND2_X1 port map( A1 => n3249, A2 => n3587, ZN => n3251);
   U2915 : INV_X1 port map( A => n3245, ZN => n3248);
   U2916 : MUX2_X1 port map( A => CWP_3_port, B => ADD_RD1(3), S => n3239, Z =>
                           n3245);
   U2917 : AOI22_X1 port map( A1 => n3252, A2 => n3588, B1 => n3253, B2 => 
                           n1815, ZN => n3246);
   U2918 : AOI21_X1 port map( B1 => CWP_1_port, B2 => n3254, A => n3239, ZN => 
                           n3252);
   U2919 : INV_X1 port map( A => n3253, ZN => n3254);
   U2920 : NOR2_X1 port map( A1 => n3237, A2 => CWP_0_port, ZN => n3253);
   U2921 : NAND2_X1 port map( A1 => n3589, A2 => n3244, ZN => n3237);
   U2922 : NOR2_X1 port map( A1 => n3249, A2 => n3587, ZN => n3226);
   U2923 : MUX2_X1 port map( A => n1814, B => n3255, S => n3239, Z => n3249);
   U2924 : INV_X1 port map( A => ADD_RD1(2), ZN => n3255);
   U2925 : NAND3_X1 port map( A1 => CWP_4_port, A2 => n2080, A3 => n3244, ZN =>
                           n3223);
   U2926 : INV_X1 port map( A => n3238, ZN => n3242);
   U2927 : AOI22_X1 port map( A1 => n3256, A2 => n3585, B1 => n3584, B2 => 
                           n3257, ZN => n3240);
   U2928 : NOR2_X1 port map( A1 => n3238, A2 => CWP_4_port, ZN => n3256);
   U2929 : NOR2_X1 port map( A1 => n3257, A2 => n3584, ZN => n3238);
   U2930 : NAND2_X1 port map( A1 => n3244, A2 => n2239, ZN => n3257);
   U2931 : OAI21_X1 port map( B1 => n1258, B2 => n2377, A => n2378, ZN => n1425
                           );
   U2932 : NAND3_X1 port map( A1 => n2377, A2 => n2374, A3 => n2389, ZN => 
                           n2378);
   U2933 : NAND2_X1 port map( A1 => n3066, A2 => n3258, ZN => n2377);
   U2934 : OAI21_X1 port map( B1 => n3259, B2 => n2222, A => n2466, ZN => n3258
                           );
   U2935 : NOR2_X1 port map( A1 => n2400, A2 => U3_U20_Z_0, ZN => n2466);
   U2936 : NAND2_X1 port map( A1 => ENABLE, A2 => n3260, ZN => n2400);
   U2937 : NOR3_X1 port map( A1 => CWP_3_port, A2 => n1812, A3 => n2375, ZN => 
                           n3259);
   U2938 : NAND4_X1 port map( A1 => n3590, A2 => n1814, A3 => n1816, A4 => 
                           n1815, ZN => n2375);
   U2939 : OAI21_X1 port map( B1 => RESET, B2 => n3261, A => n3065, ZN => n3066
                           );
   U2940 : OAI21_X1 port map( B1 => n3583, B2 => n2390, A => n2374, ZN => n3065
                           );
   U2941 : INV_X1 port map( A => ENABLE, ZN => n2390);
   U2942 : NOR2_X1 port map( A1 => n1812, A2 => U3_U4_Z_0, ZN => U3_U3_Z_5);
   U2943 : NAND2_X1 port map( A1 => n1813, A2 => n2526, ZN => U3_U3_Z_3);
   U2944 : NAND2_X1 port map( A1 => n1814, A2 => n2526, ZN => U3_U3_Z_2);
   U2945 : NOR2_X1 port map( A1 => n1815, A2 => U3_U4_Z_0, ZN => U3_U3_Z_1);
   U2946 : NOR2_X1 port map( A1 => n1816, A2 => U3_U4_Z_0, ZN => U3_U3_Z_0);
   U2947 : INV_X1 port map( A => n2526, ZN => U3_U4_Z_0);
   U2948 : NAND2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), ZN => n2526);
   U2949 : OR2_X1 port map( A1 => n3262, A2 => n3263, ZN => U3_U23_Z_0);
   U2950 : OAI21_X1 port map( B1 => n3264, B2 => n2992, A => n3265, ZN => 
                           U3_U22_Z_3);
   U2951 : INV_X1 port map( A => ADD_RD2(3), ZN => n2992);
   U2952 : NOR2_X1 port map( A1 => n3025, A2 => n2991, ZN => U3_U22_Z_2);
   U2953 : INV_X1 port map( A => ADD_RD2(2), ZN => n2991);
   U2954 : NOR2_X1 port map( A1 => n3025, A2 => n3022, ZN => U3_U22_Z_1);
   U2955 : INV_X1 port map( A => ADD_RD2(1), ZN => n3022);
   U2956 : OAI21_X1 port map( B1 => n3025, B2 => n3021, A => n3266, ZN => 
                           U3_U22_Z_0);
   U2957 : INV_X1 port map( A => ADD_RD2(0), ZN => n3021);
   U2958 : NAND3_X1 port map( A1 => n3267, A2 => n3268, A3 => n3269, ZN => 
                           U3_U21_Z_5);
   U2959 : AOI22_X1 port map( A1 => n3263, A2 => n3584, B1 => n3262, B2 => 
                           n2239, ZN => n3269);
   U2960 : NAND3_X1 port map( A1 => n2387, A2 => n2189, A3 => n3585, ZN => 
                           n3268);
   U2961 : OAI21_X1 port map( B1 => n3270, B2 => n3271, A => CWP_4_port, ZN => 
                           n3267);
   U2962 : OAI22_X1 port map( A1 => n1812, A2 => n3272, B1 => n3266, B2 => 
                           n2080, ZN => U3_U21_Z_4);
   U2963 : OAI22_X1 port map( A1 => n1813, A2 => n3272, B1 => n3266, B2 => 
                           n2081, ZN => U3_U21_Z_3);
   U2964 : OAI22_X1 port map( A1 => n1814, A2 => n3272, B1 => n3266, B2 => 
                           n2187, ZN => U3_U21_Z_2);
   U2965 : OAI22_X1 port map( A1 => n1815, A2 => n3272, B1 => n3266, B2 => 
                           n2082, ZN => U3_U21_Z_1);
   U2966 : OAI22_X1 port map( A1 => n1816, A2 => n3272, B1 => n3266, B2 => 
                           n2188, ZN => U3_U21_Z_0);
   U2967 : AOI21_X1 port map( B1 => n2387, B2 => n2189, A => n3263, ZN => n3266
                           );
   U2968 : NOR2_X1 port map( A1 => n3273, A2 => n2392, ZN => n3263);
   U2969 : NOR3_X1 port map( A1 => n2557, A2 => n3584, A3 => n2486, ZN => n2392
                           );
   U2970 : NAND3_X1 port map( A1 => n2081, A2 => n2080, A3 => n2187, ZN => 
                           n2486);
   U2971 : INV_X1 port map( A => n2570, ZN => n3273);
   U2972 : NOR3_X1 port map( A1 => n3261, A2 => n3582, A3 => n2189, ZN => n2570
                           );
   U2973 : INV_X1 port map( A => n2387, ZN => n3261);
   U2974 : NAND3_X1 port map( A1 => n3274, A2 => n2187, A3 => n3581, ZN => 
                           n2387);
   U2975 : INV_X1 port map( A => n2557, ZN => n3274);
   U2976 : NAND2_X1 port map( A1 => n2082, A2 => n2188, ZN => n2557);
   U2977 : NOR3_X1 port map( A1 => n3262, A2 => n3271, A3 => n3270, ZN => n3272
                           );
   U2978 : NOR2_X1 port map( A1 => n3265, A2 => U3_U20_Z_0, ZN => n3270);
   U2979 : INV_X1 port map( A => n3025, ZN => n3271);
   U2980 : NAND2_X1 port map( A1 => n3239, A2 => n2389, ZN => n3025);
   U2981 : AND2_X1 port map( A1 => n3260, A2 => U3_U20_Z_0, ZN => n3262);
   U2982 : INV_X1 port map( A => n3265, ZN => n3260);
   U2983 : NAND2_X1 port map( A1 => n2389, A2 => n3244, ZN => n3265);
   U2984 : INV_X1 port map( A => n3239, ZN => n3244);
   U2985 : NOR2_X1 port map( A1 => RET, A2 => CALL, ZN => n3239);
   U2986 : INV_X1 port map( A => n3264, ZN => n2389);
   U2987 : NAND2_X1 port map( A1 => n3582, A2 => n3583, ZN => n3264);
   U2988 : INV_X1 port map( A => RET, ZN => n3275);

end SYN_Behavioral;
